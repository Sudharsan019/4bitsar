VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_4Bit_SAR_ADC
  CLASS BLOCK ;
  FOREIGN tt_um_4Bit_SAR_ADC ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.000000 ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.000000 ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 90.995 197.375 91.165 197.565 ;
        RECT 93.285 197.375 93.455 197.565 ;
        RECT 94.665 197.375 94.835 197.565 ;
        RECT 95.130 197.425 95.250 197.535 ;
        RECT 95.595 197.375 95.765 197.565 ;
        RECT 97.435 197.375 97.605 197.565 ;
        RECT 102.965 197.420 103.125 197.530 ;
        RECT 104.335 197.375 104.505 197.565 ;
        RECT 109.855 197.375 110.025 197.565 ;
        RECT 115.375 197.375 115.545 197.565 ;
        RECT 117.215 197.375 117.385 197.565 ;
        RECT 119.975 197.375 120.145 197.565 ;
        RECT 90.855 196.565 92.225 197.375 ;
        RECT 92.235 196.595 93.605 197.375 ;
        RECT 93.615 196.595 94.985 197.375 ;
        RECT 95.455 196.695 97.285 197.375 ;
        RECT 95.940 196.465 97.285 196.695 ;
        RECT 97.295 196.565 102.805 197.375 ;
        RECT 103.745 196.505 104.175 197.290 ;
        RECT 104.195 196.565 109.705 197.375 ;
        RECT 109.715 196.565 115.225 197.375 ;
        RECT 115.235 196.565 116.605 197.375 ;
        RECT 116.625 196.505 117.055 197.290 ;
        RECT 117.075 196.565 118.905 197.375 ;
        RECT 118.915 196.565 120.285 197.375 ;
      LAYER nwell ;
        RECT 90.660 193.345 120.480 196.175 ;
      LAYER pwell ;
        RECT 90.855 192.145 92.225 192.955 ;
        RECT 92.235 192.145 97.745 192.955 ;
        RECT 97.755 192.145 103.265 192.955 ;
        RECT 103.745 192.230 104.175 193.015 ;
        RECT 104.195 192.145 109.705 192.955 ;
        RECT 109.715 192.145 118.820 192.825 ;
        RECT 118.915 192.145 120.285 192.955 ;
        RECT 90.995 191.935 91.165 192.145 ;
        RECT 92.375 191.935 92.545 192.145 ;
        RECT 97.895 192.125 98.065 192.145 ;
        RECT 97.895 191.955 98.070 192.125 ;
        RECT 103.410 191.985 103.530 192.095 ;
        RECT 104.335 191.955 104.505 192.145 ;
        RECT 97.900 191.935 98.070 191.955 ;
        RECT 109.855 191.935 110.025 192.145 ;
        RECT 115.375 191.935 115.545 192.125 ;
        RECT 117.215 191.935 117.385 192.125 ;
        RECT 119.975 191.935 120.145 192.145 ;
        RECT 90.855 191.125 92.225 191.935 ;
        RECT 92.235 191.125 97.745 191.935 ;
        RECT 97.755 191.255 109.705 191.935 ;
        RECT 101.660 191.035 103.930 191.255 ;
        RECT 105.535 191.035 109.705 191.255 ;
        RECT 109.715 191.125 115.225 191.935 ;
        RECT 115.235 191.125 116.605 191.935 ;
        RECT 116.625 191.065 117.055 191.850 ;
        RECT 117.075 191.125 118.905 191.935 ;
        RECT 118.915 191.125 120.285 191.935 ;
        RECT 107.370 191.025 109.705 191.035 ;
      LAYER nwell ;
        RECT 90.660 187.905 120.480 190.735 ;
      LAYER pwell ;
        RECT 90.855 186.705 92.225 187.515 ;
        RECT 97.665 187.385 98.595 187.605 ;
        RECT 101.315 187.385 103.670 187.615 ;
        RECT 93.155 186.705 103.670 187.385 ;
        RECT 103.745 186.790 104.175 187.575 ;
        RECT 104.250 187.385 106.605 187.615 ;
        RECT 109.325 187.385 110.255 187.605 ;
        RECT 104.250 186.705 114.765 187.385 ;
        RECT 114.775 186.705 118.445 187.515 ;
        RECT 118.915 186.705 120.285 187.515 ;
        RECT 90.995 186.495 91.165 186.705 ;
        RECT 93.295 186.685 93.465 186.705 ;
        RECT 92.385 186.550 92.545 186.660 ;
        RECT 93.285 186.515 93.465 186.685 ;
        RECT 93.285 186.495 93.455 186.515 ;
        RECT 93.755 186.495 93.925 186.685 ;
        RECT 99.275 186.495 99.445 186.685 ;
        RECT 112.610 186.495 112.780 186.685 ;
        RECT 113.075 186.495 113.245 186.685 ;
        RECT 114.455 186.515 114.625 186.705 ;
        RECT 114.915 186.515 115.085 186.705 ;
        RECT 117.210 186.545 117.330 186.655 ;
        RECT 118.585 186.495 118.755 186.685 ;
        RECT 119.975 186.495 120.145 186.705 ;
        RECT 90.855 185.685 92.225 186.495 ;
        RECT 92.235 185.715 93.605 186.495 ;
        RECT 93.615 185.685 99.125 186.495 ;
        RECT 99.135 185.685 100.965 186.495 ;
        RECT 100.975 185.815 112.925 186.495 ;
        RECT 100.975 185.595 105.145 185.815 ;
        RECT 106.750 185.595 109.020 185.815 ;
        RECT 112.935 185.685 116.605 186.495 ;
        RECT 116.625 185.625 117.055 186.410 ;
        RECT 117.535 185.715 118.905 186.495 ;
        RECT 118.915 185.685 120.285 186.495 ;
        RECT 100.975 185.585 103.310 185.595 ;
      LAYER nwell ;
        RECT 90.660 182.465 120.480 185.295 ;
      LAYER pwell ;
        RECT 90.855 181.265 92.225 182.075 ;
        RECT 97.665 181.945 98.595 182.165 ;
        RECT 101.315 181.945 103.670 182.175 ;
        RECT 104.195 182.165 106.530 182.175 ;
        RECT 93.155 181.265 103.670 181.945 ;
        RECT 103.745 181.350 104.175 182.135 ;
        RECT 104.195 181.945 108.365 182.165 ;
        RECT 109.970 181.945 112.240 182.165 ;
        RECT 104.195 181.265 116.145 181.945 ;
        RECT 116.155 181.265 118.905 182.075 ;
        RECT 118.915 181.265 120.285 182.075 ;
        RECT 90.995 181.055 91.165 181.265 ;
        RECT 92.375 181.055 92.545 181.245 ;
        RECT 93.295 181.075 93.465 181.265 ;
        RECT 96.065 181.100 96.225 181.210 ;
        RECT 108.470 181.055 108.640 181.245 ;
        RECT 108.935 181.055 109.105 181.245 ;
        RECT 114.455 181.055 114.625 181.245 ;
        RECT 115.830 181.075 116.000 181.265 ;
        RECT 116.295 181.215 116.465 181.265 ;
        RECT 116.290 181.105 116.465 181.215 ;
        RECT 116.295 181.075 116.465 181.105 ;
        RECT 117.215 181.055 117.385 181.245 ;
        RECT 119.975 181.055 120.145 181.265 ;
        RECT 90.855 180.245 92.225 181.055 ;
        RECT 92.235 180.245 95.905 181.055 ;
        RECT 96.835 180.375 108.785 181.055 ;
        RECT 96.835 180.155 101.005 180.375 ;
        RECT 102.610 180.155 104.880 180.375 ;
        RECT 108.795 180.245 114.305 181.055 ;
        RECT 114.315 180.245 116.145 181.055 ;
        RECT 116.625 180.185 117.055 180.970 ;
        RECT 117.075 180.245 118.905 181.055 ;
        RECT 118.915 180.245 120.285 181.055 ;
        RECT 96.835 180.145 99.170 180.155 ;
      LAYER nwell ;
        RECT 90.660 177.025 120.480 179.855 ;
      LAYER pwell ;
        RECT 90.855 175.825 92.225 176.635 ;
        RECT 97.665 176.505 98.595 176.725 ;
        RECT 101.315 176.505 103.670 176.735 ;
        RECT 93.155 175.825 103.670 176.505 ;
        RECT 103.745 175.910 104.175 176.695 ;
        RECT 104.565 176.625 106.910 176.735 ;
        RECT 104.565 176.505 107.840 176.625 ;
        RECT 112.485 176.505 113.405 176.725 ;
        RECT 104.565 175.825 114.765 176.505 ;
        RECT 114.775 175.825 118.445 176.635 ;
        RECT 118.915 175.825 120.285 176.635 ;
        RECT 90.995 175.615 91.165 175.825 ;
        RECT 93.295 175.805 93.465 175.825 ;
        RECT 92.385 175.670 92.545 175.780 ;
        RECT 93.285 175.635 93.465 175.805 ;
        RECT 93.285 175.615 93.455 175.635 ;
        RECT 94.665 175.615 94.835 175.805 ;
        RECT 95.145 175.660 95.305 175.770 ;
        RECT 107.550 175.615 107.720 175.805 ;
        RECT 108.015 175.615 108.185 175.805 ;
        RECT 113.535 175.615 113.705 175.805 ;
        RECT 114.455 175.635 114.625 175.825 ;
        RECT 114.915 175.635 115.085 175.825 ;
        RECT 116.290 175.665 116.410 175.775 ;
        RECT 117.215 175.615 117.385 175.805 ;
        RECT 118.590 175.665 118.710 175.775 ;
        RECT 119.975 175.615 120.145 175.825 ;
        RECT 90.855 174.805 92.225 175.615 ;
        RECT 92.235 174.835 93.605 175.615 ;
        RECT 93.615 174.835 94.985 175.615 ;
        RECT 95.915 174.935 107.865 175.615 ;
        RECT 95.915 174.715 100.085 174.935 ;
        RECT 101.690 174.715 103.960 174.935 ;
        RECT 107.875 174.805 113.385 175.615 ;
        RECT 113.395 174.805 116.145 175.615 ;
        RECT 116.625 174.745 117.055 175.530 ;
        RECT 117.075 174.805 118.905 175.615 ;
        RECT 118.915 174.805 120.285 175.615 ;
        RECT 95.915 174.705 98.250 174.715 ;
      LAYER nwell ;
        RECT 90.660 171.585 120.480 174.415 ;
      LAYER pwell ;
        RECT 90.855 170.385 92.225 171.195 ;
        RECT 92.320 170.385 101.425 171.065 ;
        RECT 102.355 170.385 103.725 171.165 ;
        RECT 103.745 170.470 104.175 171.255 ;
        RECT 104.280 170.385 113.385 171.065 ;
        RECT 113.395 170.385 116.145 171.195 ;
        RECT 116.625 170.470 117.055 171.255 ;
        RECT 117.075 170.385 118.905 171.195 ;
        RECT 118.915 170.385 120.285 171.195 ;
        RECT 90.995 170.195 91.165 170.385 ;
        RECT 101.115 170.195 101.285 170.385 ;
        RECT 101.585 170.230 101.745 170.340 ;
        RECT 103.405 170.195 103.575 170.385 ;
        RECT 113.075 170.195 113.245 170.385 ;
        RECT 113.535 170.195 113.705 170.385 ;
        RECT 116.290 170.225 116.410 170.335 ;
        RECT 117.215 170.195 117.385 170.385 ;
        RECT 119.975 170.195 120.145 170.385 ;
        RECT 48.665 146.725 52.765 153.195 ;
      LAYER nwell ;
        RECT 53.905 145.145 58.095 153.195 ;
      LAYER pwell ;
        RECT 62.195 146.700 66.295 153.170 ;
      LAYER nwell ;
        RECT 67.435 145.120 71.625 153.170 ;
      LAYER pwell ;
        RECT 76.000 146.700 80.100 153.170 ;
      LAYER nwell ;
        RECT 81.240 145.120 85.430 153.170 ;
      LAYER pwell ;
        RECT 89.690 146.700 93.790 153.170 ;
      LAYER nwell ;
        RECT 94.930 145.120 99.120 153.170 ;
      LAYER pwell ;
        RECT 66.405 137.115 68.415 138.915 ;
        RECT 66.405 136.715 70.420 137.115 ;
        RECT 74.440 136.715 76.450 136.915 ;
        RECT 66.405 121.095 76.450 136.715 ;
        RECT 87.085 130.595 98.475 136.695 ;
        RECT 99.995 130.760 107.665 136.720 ;
        RECT 109.905 132.000 112.365 134.710 ;
      LAYER nwell ;
        RECT 87.090 122.000 94.480 128.190 ;
        RECT 96.135 121.995 108.105 128.185 ;
        RECT 109.880 124.490 112.340 127.180 ;
        RECT 119.355 121.980 122.315 124.980 ;
      LAYER pwell ;
        RECT 68.410 110.475 74.440 121.095 ;
      LAYER nwell ;
        RECT 119.355 118.790 125.275 121.980 ;
        RECT 82.220 108.310 86.180 114.500 ;
        RECT 89.170 108.310 94.560 114.500 ;
        RECT 97.560 108.315 101.520 114.505 ;
      LAYER pwell ;
        RECT 119.350 114.380 125.270 117.480 ;
      LAYER nwell ;
        RECT 103.810 108.830 106.270 111.520 ;
      LAYER pwell ;
        RECT 119.350 111.380 122.310 114.380 ;
        RECT 79.930 105.650 86.180 107.650 ;
        RECT 97.560 105.650 106.270 107.645 ;
        RECT 79.930 103.745 106.270 105.650 ;
        RECT 79.930 101.550 103.810 103.745 ;
        RECT 97.560 101.545 103.810 101.550 ;
      LAYER li1 ;
        RECT 90.850 197.395 120.290 197.565 ;
        RECT 90.935 196.645 92.145 197.395 ;
        RECT 92.315 196.720 92.575 197.225 ;
        RECT 92.755 197.015 93.085 197.395 ;
        RECT 93.265 196.845 93.435 197.225 ;
        RECT 90.935 196.105 91.455 196.645 ;
        RECT 91.625 195.935 92.145 196.475 ;
        RECT 90.935 194.845 92.145 195.935 ;
        RECT 92.315 195.920 92.495 196.720 ;
        RECT 92.770 196.675 93.435 196.845 ;
        RECT 93.695 196.720 93.955 197.225 ;
        RECT 94.135 197.015 94.465 197.395 ;
        RECT 94.645 196.845 94.815 197.225 ;
        RECT 92.770 196.420 92.940 196.675 ;
        RECT 92.665 196.090 92.940 196.420 ;
        RECT 93.165 196.125 93.505 196.495 ;
        RECT 92.770 195.945 92.940 196.090 ;
        RECT 92.315 195.015 92.585 195.920 ;
        RECT 92.770 195.775 93.445 195.945 ;
        RECT 92.755 194.845 93.085 195.605 ;
        RECT 93.265 195.015 93.445 195.775 ;
        RECT 93.695 195.920 93.875 196.720 ;
        RECT 94.150 196.675 94.815 196.845 ;
        RECT 95.625 196.845 95.795 197.225 ;
        RECT 96.010 197.015 96.340 197.395 ;
        RECT 95.625 196.675 96.340 196.845 ;
        RECT 94.150 196.420 94.320 196.675 ;
        RECT 94.045 196.090 94.320 196.420 ;
        RECT 94.545 196.125 94.885 196.495 ;
        RECT 95.535 196.125 95.890 196.495 ;
        RECT 96.170 196.485 96.340 196.675 ;
        RECT 96.510 196.650 96.765 197.225 ;
        RECT 96.170 196.155 96.425 196.485 ;
        RECT 94.150 195.945 94.320 196.090 ;
        RECT 96.170 195.945 96.340 196.155 ;
        RECT 93.695 195.015 93.965 195.920 ;
        RECT 94.150 195.775 94.825 195.945 ;
        RECT 94.135 194.845 94.465 195.605 ;
        RECT 94.645 195.015 94.825 195.775 ;
        RECT 95.625 195.775 96.340 195.945 ;
        RECT 96.595 195.920 96.765 196.650 ;
        RECT 96.940 196.555 97.200 197.395 ;
        RECT 97.375 196.850 102.720 197.395 ;
        RECT 98.960 196.020 99.300 196.850 ;
        RECT 103.815 196.670 104.105 197.395 ;
        RECT 104.275 196.850 109.620 197.395 ;
        RECT 109.795 196.850 115.140 197.395 ;
        RECT 95.625 195.015 95.795 195.775 ;
        RECT 96.010 194.845 96.340 195.605 ;
        RECT 96.510 195.015 96.765 195.920 ;
        RECT 96.940 194.845 97.200 195.995 ;
        RECT 100.780 195.280 101.130 196.530 ;
        RECT 105.860 196.020 106.200 196.850 ;
        RECT 97.375 194.845 102.720 195.280 ;
        RECT 103.815 194.845 104.105 196.010 ;
        RECT 107.680 195.280 108.030 196.530 ;
        RECT 111.380 196.020 111.720 196.850 ;
        RECT 115.315 196.645 116.525 197.395 ;
        RECT 116.695 196.670 116.985 197.395 ;
        RECT 113.200 195.280 113.550 196.530 ;
        RECT 115.315 196.105 115.835 196.645 ;
        RECT 117.155 196.625 118.825 197.395 ;
        RECT 118.995 196.645 120.205 197.395 ;
        RECT 116.005 195.935 116.525 196.475 ;
        RECT 117.155 196.105 117.905 196.625 ;
        RECT 104.275 194.845 109.620 195.280 ;
        RECT 109.795 194.845 115.140 195.280 ;
        RECT 115.315 194.845 116.525 195.935 ;
        RECT 116.695 194.845 116.985 196.010 ;
        RECT 118.075 195.935 118.825 196.455 ;
        RECT 117.155 194.845 118.825 195.935 ;
        RECT 118.995 195.935 119.515 196.475 ;
        RECT 119.685 196.105 120.205 196.645 ;
        RECT 118.995 194.845 120.205 195.935 ;
        RECT 90.850 194.675 120.290 194.845 ;
        RECT 90.935 193.585 92.145 194.675 ;
        RECT 92.315 194.240 97.660 194.675 ;
        RECT 97.835 194.240 103.180 194.675 ;
        RECT 90.935 192.875 91.455 193.415 ;
        RECT 91.625 193.045 92.145 193.585 ;
        RECT 90.935 192.125 92.145 192.875 ;
        RECT 93.900 192.670 94.240 193.500 ;
        RECT 95.720 192.990 96.070 194.240 ;
        RECT 99.420 192.670 99.760 193.500 ;
        RECT 101.240 192.990 101.590 194.240 ;
        RECT 103.815 193.510 104.105 194.675 ;
        RECT 104.275 194.240 109.620 194.675 ;
        RECT 92.315 192.125 97.660 192.670 ;
        RECT 97.835 192.125 103.180 192.670 ;
        RECT 103.815 192.125 104.105 192.850 ;
        RECT 105.860 192.670 106.200 193.500 ;
        RECT 107.680 192.990 108.030 194.240 ;
        RECT 109.805 193.865 110.100 194.675 ;
        RECT 110.280 193.365 110.525 194.505 ;
        RECT 110.700 193.865 110.960 194.675 ;
        RECT 111.560 194.670 117.835 194.675 ;
        RECT 111.140 193.365 111.390 194.500 ;
        RECT 111.560 193.875 111.820 194.670 ;
        RECT 111.990 193.775 112.250 194.500 ;
        RECT 112.420 193.945 112.680 194.670 ;
        RECT 112.850 193.775 113.110 194.500 ;
        RECT 113.280 193.945 113.540 194.670 ;
        RECT 113.710 193.775 113.970 194.500 ;
        RECT 114.140 193.945 114.400 194.670 ;
        RECT 114.570 193.775 114.830 194.500 ;
        RECT 115.000 193.945 115.245 194.670 ;
        RECT 115.415 193.775 115.675 194.500 ;
        RECT 115.860 193.945 116.105 194.670 ;
        RECT 116.275 193.775 116.535 194.500 ;
        RECT 116.720 193.945 116.965 194.670 ;
        RECT 117.135 193.775 117.395 194.500 ;
        RECT 117.580 193.945 117.835 194.670 ;
        RECT 111.990 193.760 117.395 193.775 ;
        RECT 118.005 193.760 118.295 194.500 ;
        RECT 118.465 193.930 118.735 194.675 ;
        RECT 111.990 193.535 118.735 193.760 ;
        RECT 109.795 192.805 110.110 193.365 ;
        RECT 110.280 193.115 117.400 193.365 ;
        RECT 104.275 192.125 109.620 192.670 ;
        RECT 109.795 192.125 110.100 192.635 ;
        RECT 110.280 192.305 110.530 193.115 ;
        RECT 110.700 192.125 110.960 192.650 ;
        RECT 111.140 192.305 111.390 193.115 ;
        RECT 117.570 192.945 118.735 193.535 ;
        RECT 118.995 193.585 120.205 194.675 ;
        RECT 118.995 193.045 119.515 193.585 ;
        RECT 111.990 192.775 118.735 192.945 ;
        RECT 119.685 192.875 120.205 193.415 ;
        RECT 111.560 192.125 111.820 192.685 ;
        RECT 111.990 192.320 112.250 192.775 ;
        RECT 112.420 192.125 112.680 192.605 ;
        RECT 112.850 192.320 113.110 192.775 ;
        RECT 113.280 192.125 113.540 192.605 ;
        RECT 113.710 192.320 113.970 192.775 ;
        RECT 114.140 192.125 114.385 192.605 ;
        RECT 114.555 192.320 114.830 192.775 ;
        RECT 115.000 192.125 115.245 192.605 ;
        RECT 115.415 192.320 115.675 192.775 ;
        RECT 115.855 192.125 116.105 192.605 ;
        RECT 116.275 192.320 116.535 192.775 ;
        RECT 116.715 192.125 116.965 192.605 ;
        RECT 117.135 192.320 117.395 192.775 ;
        RECT 117.575 192.125 117.835 192.605 ;
        RECT 118.005 192.320 118.265 192.775 ;
        RECT 118.435 192.125 118.735 192.605 ;
        RECT 118.995 192.125 120.205 192.875 ;
        RECT 90.850 191.955 120.290 192.125 ;
        RECT 90.935 191.205 92.145 191.955 ;
        RECT 92.315 191.410 97.660 191.955 ;
        RECT 90.935 190.665 91.455 191.205 ;
        RECT 91.625 190.495 92.145 191.035 ;
        RECT 93.900 190.580 94.240 191.410 ;
        RECT 97.835 191.405 98.095 191.695 ;
        RECT 98.265 191.575 98.595 191.955 ;
        RECT 97.835 191.235 98.590 191.405 ;
        RECT 90.935 189.405 92.145 190.495 ;
        RECT 95.720 189.840 96.070 191.090 ;
        RECT 97.835 190.415 98.190 191.065 ;
        RECT 98.360 190.245 98.590 191.235 ;
        RECT 97.835 190.075 98.590 190.245 ;
        RECT 92.315 189.405 97.660 189.840 ;
        RECT 97.835 189.575 98.095 190.075 ;
        RECT 98.265 189.405 98.595 189.905 ;
        RECT 98.765 189.575 98.990 191.695 ;
        RECT 99.185 191.575 99.535 191.955 ;
        RECT 99.705 191.405 99.875 191.735 ;
        RECT 100.155 191.575 101.150 191.775 ;
        RECT 99.160 191.215 99.875 191.405 ;
        RECT 99.160 190.245 99.330 191.215 ;
        RECT 99.500 190.415 99.910 191.035 ;
        RECT 100.080 190.465 100.300 191.335 ;
        RECT 100.480 191.025 100.810 191.395 ;
        RECT 100.980 190.845 101.150 191.575 ;
        RECT 101.320 191.515 101.490 191.955 ;
        RECT 101.660 191.615 102.830 191.785 ;
        RECT 101.660 191.495 101.990 191.615 ;
        RECT 101.340 191.075 101.750 191.305 ;
        RECT 102.160 191.275 102.490 191.445 ;
        RECT 102.660 191.325 102.830 191.615 ;
        RECT 103.100 191.575 103.430 191.955 ;
        RECT 104.070 191.575 104.835 191.775 ;
        RECT 102.270 191.145 102.490 191.275 ;
        RECT 101.340 190.975 101.670 191.075 ;
        RECT 102.270 190.975 103.580 191.145 ;
        RECT 100.750 190.805 101.150 190.845 ;
        RECT 101.880 190.805 102.100 190.885 ;
        RECT 100.750 190.635 102.100 190.805 ;
        RECT 99.160 190.075 99.875 190.245 ;
        RECT 100.080 190.085 100.580 190.465 ;
        RECT 99.185 189.405 99.535 189.905 ;
        RECT 99.705 189.575 99.875 190.075 ;
        RECT 100.750 189.790 100.920 190.635 ;
        RECT 101.850 190.555 102.100 190.635 ;
        RECT 101.090 190.255 101.340 190.465 ;
        RECT 102.270 190.255 102.440 190.975 ;
        RECT 103.250 190.805 103.580 190.975 ;
        RECT 103.875 190.915 104.160 191.335 ;
        RECT 102.610 190.625 102.940 190.805 ;
        RECT 103.875 190.735 104.495 190.915 ;
        RECT 102.610 190.385 103.615 190.625 ;
        RECT 101.090 190.005 102.440 190.255 ;
        RECT 100.090 189.620 100.920 189.790 ;
        RECT 101.160 189.405 101.540 189.835 ;
        RECT 101.840 189.665 102.010 190.005 ;
        RECT 102.630 189.405 102.960 190.125 ;
        RECT 103.815 190.055 104.050 190.465 ;
        RECT 104.290 190.135 104.495 190.735 ;
        RECT 104.665 190.805 104.835 191.575 ;
        RECT 105.015 191.515 105.275 191.955 ;
        RECT 105.535 191.615 106.705 191.785 ;
        RECT 105.535 191.495 105.865 191.615 ;
        RECT 106.535 191.455 106.705 191.615 ;
        RECT 105.210 190.975 105.585 191.305 ;
        RECT 106.035 191.260 106.365 191.445 ;
        RECT 106.990 191.285 107.225 191.775 ;
        RECT 105.795 190.805 106.015 190.965 ;
        RECT 104.665 190.635 106.015 190.805 ;
        RECT 104.665 189.790 104.835 190.635 ;
        RECT 105.005 190.125 105.255 190.465 ;
        RECT 106.185 190.125 106.365 191.260 ;
        RECT 106.535 191.115 107.225 191.285 ;
        RECT 107.450 191.235 107.780 191.955 ;
        RECT 107.950 191.325 108.235 191.785 ;
        RECT 106.535 190.465 106.810 191.115 ;
        RECT 107.065 190.715 107.440 190.945 ;
        RECT 107.610 190.715 107.860 191.045 ;
        RECT 106.535 190.295 107.295 190.465 ;
        RECT 107.610 190.125 107.780 190.715 ;
        RECT 108.030 190.410 108.235 191.325 ;
        RECT 105.005 189.955 107.780 190.125 ;
        RECT 104.005 189.620 104.835 189.790 ;
        RECT 105.075 189.405 105.455 189.785 ;
        RECT 105.695 189.665 105.865 189.955 ;
        RECT 106.395 189.405 107.780 189.785 ;
        RECT 107.950 189.575 108.235 190.410 ;
        RECT 108.405 191.045 108.720 191.785 ;
        RECT 108.900 191.495 109.195 191.955 ;
        RECT 109.365 191.215 109.625 191.785 ;
        RECT 109.795 191.410 115.140 191.955 ;
        RECT 108.405 190.715 109.240 191.045 ;
        RECT 108.405 189.625 108.720 190.715 ;
        RECT 109.410 190.595 109.625 191.215 ;
        RECT 108.900 189.405 109.195 190.275 ;
        RECT 109.365 189.575 109.625 190.595 ;
        RECT 111.380 190.580 111.720 191.410 ;
        RECT 115.315 191.205 116.525 191.955 ;
        RECT 116.695 191.230 116.985 191.955 ;
        RECT 113.200 189.840 113.550 191.090 ;
        RECT 115.315 190.665 115.835 191.205 ;
        RECT 117.155 191.185 118.825 191.955 ;
        RECT 118.995 191.205 120.205 191.955 ;
        RECT 116.005 190.495 116.525 191.035 ;
        RECT 117.155 190.665 117.905 191.185 ;
        RECT 109.795 189.405 115.140 189.840 ;
        RECT 115.315 189.405 116.525 190.495 ;
        RECT 116.695 189.405 116.985 190.570 ;
        RECT 118.075 190.495 118.825 191.015 ;
        RECT 117.155 189.405 118.825 190.495 ;
        RECT 118.995 190.495 119.515 191.035 ;
        RECT 119.685 190.665 120.205 191.205 ;
        RECT 118.995 189.405 120.205 190.495 ;
        RECT 90.850 189.235 120.290 189.405 ;
        RECT 90.935 188.145 92.145 189.235 ;
        RECT 93.240 188.565 93.495 189.065 ;
        RECT 93.665 188.735 93.995 189.235 ;
        RECT 93.240 188.395 93.990 188.565 ;
        RECT 90.935 187.435 91.455 187.975 ;
        RECT 91.625 187.605 92.145 188.145 ;
        RECT 93.240 187.575 93.590 188.225 ;
        RECT 90.935 186.685 92.145 187.435 ;
        RECT 93.760 187.405 93.990 188.395 ;
        RECT 93.240 187.235 93.990 187.405 ;
        RECT 93.240 186.945 93.495 187.235 ;
        RECT 93.665 186.685 93.995 187.065 ;
        RECT 94.165 186.945 94.335 189.065 ;
        RECT 94.505 188.265 94.830 189.050 ;
        RECT 95.000 188.775 95.250 189.235 ;
        RECT 95.420 188.735 95.670 189.065 ;
        RECT 95.885 188.735 96.565 189.065 ;
        RECT 95.420 188.605 95.590 188.735 ;
        RECT 95.195 188.435 95.590 188.605 ;
        RECT 94.565 187.215 95.025 188.265 ;
        RECT 95.195 187.075 95.365 188.435 ;
        RECT 95.760 188.175 96.225 188.565 ;
        RECT 95.535 187.365 95.885 187.985 ;
        RECT 96.055 187.585 96.225 188.175 ;
        RECT 96.395 187.955 96.565 188.735 ;
        RECT 96.735 188.635 96.905 188.975 ;
        RECT 97.140 188.805 97.470 189.235 ;
        RECT 97.640 188.635 97.810 188.975 ;
        RECT 98.105 188.775 98.475 189.235 ;
        RECT 96.735 188.465 97.810 188.635 ;
        RECT 98.645 188.605 98.815 189.065 ;
        RECT 99.050 188.725 99.920 189.065 ;
        RECT 100.090 188.775 100.340 189.235 ;
        RECT 98.255 188.435 98.815 188.605 ;
        RECT 98.255 188.295 98.425 188.435 ;
        RECT 96.925 188.125 98.425 188.295 ;
        RECT 99.120 188.265 99.580 188.555 ;
        RECT 96.395 187.785 98.085 187.955 ;
        RECT 96.055 187.365 96.410 187.585 ;
        RECT 96.580 187.075 96.750 187.785 ;
        RECT 96.955 187.365 97.745 187.615 ;
        RECT 97.915 187.605 98.085 187.785 ;
        RECT 98.255 187.435 98.425 188.125 ;
        RECT 94.695 186.685 95.025 187.045 ;
        RECT 95.195 186.905 95.690 187.075 ;
        RECT 95.895 186.905 96.750 187.075 ;
        RECT 97.625 186.685 97.955 187.145 ;
        RECT 98.165 187.045 98.425 187.435 ;
        RECT 98.615 188.255 99.580 188.265 ;
        RECT 99.750 188.345 99.920 188.725 ;
        RECT 100.510 188.685 100.680 188.975 ;
        RECT 100.860 188.855 101.580 189.235 ;
        RECT 100.510 188.515 101.310 188.685 ;
        RECT 98.615 188.095 99.290 188.255 ;
        RECT 99.750 188.175 100.970 188.345 ;
        RECT 98.615 187.305 98.825 188.095 ;
        RECT 99.750 188.085 99.920 188.175 ;
        RECT 98.995 187.305 99.345 187.925 ;
        RECT 99.515 187.915 99.920 188.085 ;
        RECT 99.515 187.135 99.685 187.915 ;
        RECT 99.855 187.465 100.075 187.745 ;
        RECT 100.255 187.635 100.795 188.005 ;
        RECT 101.140 187.925 101.310 188.515 ;
        RECT 101.750 188.055 102.155 189.065 ;
        RECT 101.805 188.045 102.155 188.055 ;
        RECT 101.140 187.895 101.585 187.925 ;
        RECT 99.855 187.295 100.385 187.465 ;
        RECT 98.165 186.875 98.515 187.045 ;
        RECT 98.735 186.855 99.685 187.135 ;
        RECT 99.855 186.685 100.045 187.125 ;
        RECT 100.215 187.065 100.385 187.295 ;
        RECT 100.555 187.235 100.795 187.635 ;
        RECT 100.965 187.595 101.585 187.895 ;
        RECT 100.965 187.420 101.290 187.595 ;
        RECT 100.965 187.065 101.285 187.420 ;
        RECT 100.215 186.895 101.285 187.065 ;
        RECT 101.485 186.685 101.655 187.370 ;
        RECT 101.825 186.875 102.155 188.045 ;
        RECT 102.345 187.925 102.675 189.025 ;
        RECT 102.910 188.095 103.080 189.235 ;
        RECT 103.330 188.045 103.585 188.925 ;
        RECT 103.815 188.070 104.105 189.235 ;
        RECT 102.345 187.595 103.205 187.925 ;
        RECT 102.345 186.945 102.595 187.595 ;
        RECT 103.375 187.395 103.585 188.045 ;
        RECT 104.335 188.045 104.590 188.925 ;
        RECT 104.840 188.095 105.010 189.235 ;
        RECT 102.910 186.685 103.080 187.280 ;
        RECT 103.330 186.865 103.585 187.395 ;
        RECT 103.815 186.685 104.105 187.410 ;
        RECT 104.335 187.395 104.545 188.045 ;
        RECT 105.245 187.925 105.575 189.025 ;
        RECT 104.715 187.595 105.575 187.925 ;
        RECT 104.335 186.865 104.590 187.395 ;
        RECT 104.840 186.685 105.010 187.280 ;
        RECT 105.325 186.945 105.575 187.595 ;
        RECT 105.765 188.055 106.170 189.065 ;
        RECT 106.340 188.855 107.060 189.235 ;
        RECT 107.240 188.685 107.410 188.975 ;
        RECT 107.580 188.775 107.830 189.235 ;
        RECT 106.610 188.515 107.410 188.685 ;
        RECT 108.000 188.725 108.870 189.065 ;
        RECT 105.765 186.875 106.095 188.055 ;
        RECT 106.610 187.925 106.780 188.515 ;
        RECT 108.000 188.345 108.170 188.725 ;
        RECT 109.105 188.605 109.275 189.065 ;
        RECT 109.445 188.775 109.815 189.235 ;
        RECT 110.110 188.635 110.280 188.975 ;
        RECT 110.450 188.805 110.780 189.235 ;
        RECT 111.015 188.635 111.185 188.975 ;
        RECT 106.950 188.175 108.170 188.345 ;
        RECT 108.340 188.265 108.800 188.555 ;
        RECT 109.105 188.435 109.665 188.605 ;
        RECT 110.110 188.465 111.185 188.635 ;
        RECT 111.355 188.735 112.035 189.065 ;
        RECT 112.250 188.735 112.500 189.065 ;
        RECT 112.670 188.775 112.920 189.235 ;
        RECT 109.495 188.295 109.665 188.435 ;
        RECT 108.340 188.255 109.305 188.265 ;
        RECT 108.000 188.085 108.170 188.175 ;
        RECT 108.630 188.095 109.305 188.255 ;
        RECT 106.335 187.895 106.780 187.925 ;
        RECT 106.335 187.595 106.955 187.895 ;
        RECT 106.630 187.420 106.955 187.595 ;
        RECT 106.265 186.685 106.435 187.370 ;
        RECT 106.635 187.065 106.955 187.420 ;
        RECT 107.125 187.635 107.665 188.005 ;
        RECT 108.000 187.915 108.405 188.085 ;
        RECT 107.125 187.235 107.365 187.635 ;
        RECT 107.845 187.465 108.065 187.745 ;
        RECT 107.535 187.295 108.065 187.465 ;
        RECT 107.535 187.065 107.705 187.295 ;
        RECT 108.235 187.135 108.405 187.915 ;
        RECT 108.575 187.305 108.925 187.925 ;
        RECT 109.095 187.305 109.305 188.095 ;
        RECT 109.495 188.125 110.995 188.295 ;
        RECT 109.495 187.435 109.665 188.125 ;
        RECT 111.355 187.955 111.525 188.735 ;
        RECT 112.330 188.605 112.500 188.735 ;
        RECT 109.835 187.785 111.525 187.955 ;
        RECT 111.695 188.175 112.160 188.565 ;
        RECT 112.330 188.435 112.725 188.605 ;
        RECT 109.835 187.605 110.005 187.785 ;
        RECT 106.635 186.895 107.705 187.065 ;
        RECT 107.875 186.685 108.065 187.125 ;
        RECT 108.235 186.855 109.185 187.135 ;
        RECT 109.495 187.045 109.755 187.435 ;
        RECT 110.175 187.365 110.965 187.615 ;
        RECT 109.405 186.875 109.755 187.045 ;
        RECT 109.965 186.685 110.295 187.145 ;
        RECT 111.170 187.075 111.340 187.785 ;
        RECT 111.695 187.585 111.865 188.175 ;
        RECT 111.510 187.365 111.865 187.585 ;
        RECT 112.035 187.365 112.385 187.985 ;
        RECT 112.555 187.075 112.725 188.435 ;
        RECT 113.090 188.265 113.415 189.050 ;
        RECT 112.895 187.215 113.355 188.265 ;
        RECT 111.170 186.905 112.025 187.075 ;
        RECT 112.230 186.905 112.725 187.075 ;
        RECT 112.895 186.685 113.225 187.045 ;
        RECT 113.585 186.945 113.755 189.065 ;
        RECT 113.925 188.735 114.255 189.235 ;
        RECT 114.425 188.565 114.680 189.065 ;
        RECT 113.930 188.395 114.680 188.565 ;
        RECT 113.930 187.405 114.160 188.395 ;
        RECT 114.330 187.575 114.680 188.225 ;
        RECT 114.855 188.145 118.365 189.235 ;
        RECT 114.855 187.455 116.505 187.975 ;
        RECT 116.675 187.625 118.365 188.145 ;
        RECT 118.995 188.145 120.205 189.235 ;
        RECT 118.995 187.605 119.515 188.145 ;
        RECT 113.930 187.235 114.680 187.405 ;
        RECT 113.925 186.685 114.255 187.065 ;
        RECT 114.425 186.945 114.680 187.235 ;
        RECT 114.855 186.685 118.365 187.455 ;
        RECT 119.685 187.435 120.205 187.975 ;
        RECT 118.995 186.685 120.205 187.435 ;
        RECT 90.850 186.515 120.290 186.685 ;
        RECT 90.935 185.765 92.145 186.515 ;
        RECT 92.315 185.840 92.575 186.345 ;
        RECT 92.755 186.135 93.085 186.515 ;
        RECT 93.265 185.965 93.435 186.345 ;
        RECT 93.695 185.970 99.040 186.515 ;
        RECT 90.935 185.225 91.455 185.765 ;
        RECT 91.625 185.055 92.145 185.595 ;
        RECT 90.935 183.965 92.145 185.055 ;
        RECT 92.315 185.040 92.495 185.840 ;
        RECT 92.770 185.795 93.435 185.965 ;
        RECT 92.770 185.540 92.940 185.795 ;
        RECT 92.665 185.210 92.940 185.540 ;
        RECT 93.165 185.245 93.505 185.615 ;
        RECT 92.770 185.065 92.940 185.210 ;
        RECT 95.280 185.140 95.620 185.970 ;
        RECT 99.215 185.745 100.885 186.515 ;
        RECT 101.055 185.775 101.315 186.345 ;
        RECT 101.485 186.055 101.780 186.515 ;
        RECT 92.315 184.135 92.585 185.040 ;
        RECT 92.770 184.895 93.445 185.065 ;
        RECT 92.755 183.965 93.085 184.725 ;
        RECT 93.265 184.135 93.445 184.895 ;
        RECT 97.100 184.400 97.450 185.650 ;
        RECT 99.215 185.225 99.965 185.745 ;
        RECT 100.135 185.055 100.885 185.575 ;
        RECT 93.695 183.965 99.040 184.400 ;
        RECT 99.215 183.965 100.885 185.055 ;
        RECT 101.055 185.155 101.270 185.775 ;
        RECT 101.960 185.605 102.275 186.345 ;
        RECT 101.440 185.275 102.275 185.605 ;
        RECT 101.055 184.135 101.315 185.155 ;
        RECT 101.485 183.965 101.780 184.835 ;
        RECT 101.960 184.185 102.275 185.275 ;
        RECT 102.445 185.885 102.730 186.345 ;
        RECT 102.445 184.970 102.650 185.885 ;
        RECT 102.900 185.795 103.230 186.515 ;
        RECT 103.455 185.845 103.690 186.335 ;
        RECT 103.975 186.175 105.145 186.345 ;
        RECT 103.975 186.015 104.145 186.175 ;
        RECT 104.815 186.055 105.145 186.175 ;
        RECT 105.405 186.075 105.665 186.515 ;
        RECT 105.845 186.135 106.610 186.335 ;
        RECT 107.250 186.135 107.580 186.515 ;
        RECT 107.850 186.175 109.020 186.345 ;
        RECT 103.455 185.675 104.145 185.845 ;
        RECT 102.820 185.275 103.070 185.605 ;
        RECT 103.240 185.275 103.615 185.505 ;
        RECT 102.445 184.135 102.730 184.970 ;
        RECT 102.900 184.685 103.070 185.275 ;
        RECT 103.870 185.025 104.145 185.675 ;
        RECT 103.385 184.855 104.145 185.025 ;
        RECT 104.315 185.820 104.645 186.005 ;
        RECT 104.315 184.685 104.495 185.820 ;
        RECT 105.095 185.535 105.470 185.865 ;
        RECT 104.665 185.365 104.885 185.525 ;
        RECT 105.845 185.365 106.015 186.135 ;
        RECT 106.520 185.475 106.805 185.895 ;
        RECT 107.850 185.885 108.020 186.175 ;
        RECT 108.690 186.055 109.020 186.175 ;
        RECT 109.190 186.075 109.360 186.515 ;
        RECT 109.530 186.135 110.525 186.335 ;
        RECT 108.190 185.835 108.520 186.005 ;
        RECT 108.190 185.705 108.410 185.835 ;
        RECT 104.665 185.195 106.015 185.365 ;
        RECT 105.425 184.685 105.675 185.025 ;
        RECT 102.900 184.515 105.675 184.685 ;
        RECT 102.900 183.965 104.285 184.345 ;
        RECT 104.815 184.225 104.985 184.515 ;
        RECT 105.845 184.350 106.015 185.195 ;
        RECT 106.185 185.295 106.805 185.475 ;
        RECT 107.100 185.535 108.410 185.705 ;
        RECT 108.930 185.635 109.340 185.865 ;
        RECT 109.010 185.535 109.340 185.635 ;
        RECT 107.100 185.365 107.430 185.535 ;
        RECT 106.185 184.695 106.390 185.295 ;
        RECT 107.740 185.185 108.070 185.365 ;
        RECT 106.630 184.615 106.865 185.025 ;
        RECT 107.065 184.945 108.070 185.185 ;
        RECT 108.240 184.815 108.410 185.535 ;
        RECT 108.580 185.365 108.800 185.445 ;
        RECT 109.530 185.405 109.700 186.135 ;
        RECT 110.805 185.965 110.975 186.295 ;
        RECT 111.145 186.135 111.495 186.515 ;
        RECT 109.870 185.585 110.200 185.955 ;
        RECT 109.530 185.365 109.930 185.405 ;
        RECT 108.580 185.195 109.930 185.365 ;
        RECT 108.580 185.115 108.830 185.195 ;
        RECT 109.340 184.815 109.590 185.025 ;
        RECT 105.225 183.965 105.605 184.345 ;
        RECT 105.845 184.180 106.675 184.350 ;
        RECT 107.720 183.965 108.050 184.685 ;
        RECT 108.240 184.565 109.590 184.815 ;
        RECT 108.670 184.225 108.840 184.565 ;
        RECT 109.140 183.965 109.520 184.395 ;
        RECT 109.760 184.350 109.930 185.195 ;
        RECT 110.380 185.025 110.600 185.895 ;
        RECT 110.805 185.775 111.520 185.965 ;
        RECT 110.100 184.645 110.600 185.025 ;
        RECT 110.770 184.975 111.180 185.595 ;
        RECT 111.350 184.805 111.520 185.775 ;
        RECT 110.805 184.635 111.520 184.805 ;
        RECT 109.760 184.180 110.590 184.350 ;
        RECT 110.805 184.135 110.975 184.635 ;
        RECT 111.145 183.965 111.495 184.465 ;
        RECT 111.690 184.135 111.915 186.255 ;
        RECT 112.085 186.135 112.415 186.515 ;
        RECT 112.585 185.965 112.845 186.255 ;
        RECT 112.090 185.795 112.845 185.965 ;
        RECT 112.090 184.805 112.320 185.795 ;
        RECT 113.015 185.745 116.525 186.515 ;
        RECT 116.695 185.790 116.985 186.515 ;
        RECT 117.615 185.840 117.875 186.345 ;
        RECT 118.055 186.135 118.385 186.515 ;
        RECT 118.565 185.965 118.735 186.345 ;
        RECT 112.490 184.975 112.845 185.625 ;
        RECT 113.015 185.225 114.665 185.745 ;
        RECT 114.835 185.055 116.525 185.575 ;
        RECT 112.090 184.635 112.845 184.805 ;
        RECT 112.085 183.965 112.415 184.465 ;
        RECT 112.585 184.135 112.845 184.635 ;
        RECT 113.015 183.965 116.525 185.055 ;
        RECT 116.695 183.965 116.985 185.130 ;
        RECT 117.615 185.040 117.795 185.840 ;
        RECT 118.070 185.795 118.735 185.965 ;
        RECT 118.070 185.540 118.240 185.795 ;
        RECT 118.995 185.765 120.205 186.515 ;
        RECT 117.965 185.210 118.240 185.540 ;
        RECT 118.465 185.245 118.805 185.615 ;
        RECT 118.070 185.065 118.240 185.210 ;
        RECT 117.615 184.135 117.885 185.040 ;
        RECT 118.070 184.895 118.745 185.065 ;
        RECT 118.055 183.965 118.385 184.725 ;
        RECT 118.565 184.135 118.745 184.895 ;
        RECT 118.995 185.055 119.515 185.595 ;
        RECT 119.685 185.225 120.205 185.765 ;
        RECT 118.995 183.965 120.205 185.055 ;
        RECT 90.850 183.795 120.290 183.965 ;
        RECT 90.935 182.705 92.145 183.795 ;
        RECT 93.240 183.125 93.495 183.625 ;
        RECT 93.665 183.295 93.995 183.795 ;
        RECT 93.240 182.955 93.990 183.125 ;
        RECT 90.935 181.995 91.455 182.535 ;
        RECT 91.625 182.165 92.145 182.705 ;
        RECT 93.240 182.135 93.590 182.785 ;
        RECT 90.935 181.245 92.145 181.995 ;
        RECT 93.760 181.965 93.990 182.955 ;
        RECT 93.240 181.795 93.990 181.965 ;
        RECT 93.240 181.505 93.495 181.795 ;
        RECT 93.665 181.245 93.995 181.625 ;
        RECT 94.165 181.505 94.335 183.625 ;
        RECT 94.505 182.825 94.830 183.610 ;
        RECT 95.000 183.335 95.250 183.795 ;
        RECT 95.420 183.295 95.670 183.625 ;
        RECT 95.885 183.295 96.565 183.625 ;
        RECT 95.420 183.165 95.590 183.295 ;
        RECT 95.195 182.995 95.590 183.165 ;
        RECT 94.565 181.775 95.025 182.825 ;
        RECT 95.195 181.635 95.365 182.995 ;
        RECT 95.760 182.735 96.225 183.125 ;
        RECT 95.535 181.925 95.885 182.545 ;
        RECT 96.055 182.145 96.225 182.735 ;
        RECT 96.395 182.515 96.565 183.295 ;
        RECT 96.735 183.195 96.905 183.535 ;
        RECT 97.140 183.365 97.470 183.795 ;
        RECT 97.640 183.195 97.810 183.535 ;
        RECT 98.105 183.335 98.475 183.795 ;
        RECT 96.735 183.025 97.810 183.195 ;
        RECT 98.645 183.165 98.815 183.625 ;
        RECT 99.050 183.285 99.920 183.625 ;
        RECT 100.090 183.335 100.340 183.795 ;
        RECT 98.255 182.995 98.815 183.165 ;
        RECT 98.255 182.855 98.425 182.995 ;
        RECT 96.925 182.685 98.425 182.855 ;
        RECT 99.120 182.825 99.580 183.115 ;
        RECT 96.395 182.345 98.085 182.515 ;
        RECT 96.055 181.925 96.410 182.145 ;
        RECT 96.580 181.635 96.750 182.345 ;
        RECT 96.955 181.925 97.745 182.175 ;
        RECT 97.915 182.165 98.085 182.345 ;
        RECT 98.255 181.995 98.425 182.685 ;
        RECT 94.695 181.245 95.025 181.605 ;
        RECT 95.195 181.465 95.690 181.635 ;
        RECT 95.895 181.465 96.750 181.635 ;
        RECT 97.625 181.245 97.955 181.705 ;
        RECT 98.165 181.605 98.425 181.995 ;
        RECT 98.615 182.815 99.580 182.825 ;
        RECT 99.750 182.905 99.920 183.285 ;
        RECT 100.510 183.245 100.680 183.535 ;
        RECT 100.860 183.415 101.580 183.795 ;
        RECT 100.510 183.075 101.310 183.245 ;
        RECT 98.615 182.655 99.290 182.815 ;
        RECT 99.750 182.735 100.970 182.905 ;
        RECT 98.615 181.865 98.825 182.655 ;
        RECT 99.750 182.645 99.920 182.735 ;
        RECT 98.995 181.865 99.345 182.485 ;
        RECT 99.515 182.475 99.920 182.645 ;
        RECT 99.515 181.695 99.685 182.475 ;
        RECT 99.855 182.025 100.075 182.305 ;
        RECT 100.255 182.195 100.795 182.565 ;
        RECT 101.140 182.485 101.310 183.075 ;
        RECT 101.750 182.615 102.155 183.625 ;
        RECT 101.140 182.455 101.585 182.485 ;
        RECT 99.855 181.855 100.385 182.025 ;
        RECT 98.165 181.435 98.515 181.605 ;
        RECT 98.735 181.415 99.685 181.695 ;
        RECT 99.855 181.245 100.045 181.685 ;
        RECT 100.215 181.625 100.385 181.855 ;
        RECT 100.555 181.795 100.795 182.195 ;
        RECT 100.965 182.155 101.585 182.455 ;
        RECT 101.825 182.435 102.155 182.615 ;
        RECT 101.805 182.265 102.155 182.435 ;
        RECT 100.965 181.980 101.290 182.155 ;
        RECT 100.965 181.625 101.285 181.980 ;
        RECT 100.215 181.455 101.285 181.625 ;
        RECT 101.485 181.245 101.655 181.930 ;
        RECT 101.825 181.435 102.155 182.265 ;
        RECT 102.345 182.485 102.675 183.585 ;
        RECT 102.910 182.655 103.080 183.795 ;
        RECT 103.330 182.605 103.585 183.485 ;
        RECT 103.815 182.630 104.105 183.795 ;
        RECT 102.345 182.155 103.205 182.485 ;
        RECT 102.345 181.505 102.595 182.155 ;
        RECT 103.375 181.955 103.585 182.605 ;
        RECT 104.275 182.605 104.535 183.625 ;
        RECT 104.705 182.925 105.000 183.795 ;
        RECT 104.275 181.985 104.490 182.605 ;
        RECT 105.180 182.485 105.495 183.575 ;
        RECT 104.660 182.155 105.495 182.485 ;
        RECT 102.910 181.245 103.080 181.840 ;
        RECT 103.330 181.425 103.585 181.955 ;
        RECT 103.815 181.245 104.105 181.970 ;
        RECT 104.275 181.415 104.535 181.985 ;
        RECT 104.705 181.245 105.000 181.705 ;
        RECT 105.180 181.415 105.495 182.155 ;
        RECT 105.665 182.790 105.950 183.625 ;
        RECT 106.120 183.415 107.505 183.795 ;
        RECT 108.035 183.245 108.205 183.535 ;
        RECT 108.445 183.415 108.825 183.795 ;
        RECT 109.065 183.410 109.895 183.580 ;
        RECT 106.120 183.075 108.895 183.245 ;
        RECT 105.665 181.875 105.870 182.790 ;
        RECT 106.120 182.485 106.290 183.075 ;
        RECT 106.605 182.735 107.365 182.905 ;
        RECT 106.040 182.155 106.290 182.485 ;
        RECT 106.460 182.255 106.835 182.485 ;
        RECT 107.090 182.085 107.365 182.735 ;
        RECT 105.665 181.415 105.950 181.875 ;
        RECT 106.120 181.245 106.450 181.965 ;
        RECT 106.675 181.915 107.365 182.085 ;
        RECT 107.535 181.940 107.715 183.075 ;
        RECT 108.645 182.735 108.895 183.075 ;
        RECT 109.065 182.565 109.235 183.410 ;
        RECT 107.885 182.395 109.235 182.565 ;
        RECT 107.885 182.235 108.105 182.395 ;
        RECT 106.675 181.425 106.910 181.915 ;
        RECT 107.535 181.755 107.865 181.940 ;
        RECT 108.315 181.895 108.690 182.225 ;
        RECT 107.195 181.585 107.365 181.745 ;
        RECT 108.035 181.585 108.365 181.705 ;
        RECT 107.195 181.415 108.365 181.585 ;
        RECT 108.625 181.245 108.885 181.685 ;
        RECT 109.065 181.625 109.235 182.395 ;
        RECT 109.405 182.465 109.610 183.065 ;
        RECT 109.850 182.735 110.085 183.145 ;
        RECT 110.940 183.075 111.270 183.795 ;
        RECT 111.890 183.195 112.060 183.535 ;
        RECT 112.360 183.365 112.740 183.795 ;
        RECT 112.980 183.410 113.810 183.580 ;
        RECT 111.460 182.945 112.810 183.195 ;
        RECT 110.285 182.575 111.290 182.815 ;
        RECT 109.405 182.285 110.025 182.465 ;
        RECT 110.960 182.395 111.290 182.575 ;
        RECT 109.740 181.865 110.025 182.285 ;
        RECT 110.320 182.225 110.650 182.395 ;
        RECT 111.460 182.225 111.630 182.945 ;
        RECT 112.560 182.735 112.810 182.945 ;
        RECT 111.800 182.565 112.050 182.645 ;
        RECT 112.980 182.565 113.150 183.410 ;
        RECT 114.025 183.125 114.195 183.625 ;
        RECT 114.365 183.295 114.715 183.795 ;
        RECT 113.320 182.735 113.820 183.115 ;
        RECT 114.025 182.955 114.740 183.125 ;
        RECT 111.800 182.395 113.150 182.565 ;
        RECT 111.800 182.315 112.020 182.395 ;
        RECT 112.750 182.355 113.150 182.395 ;
        RECT 110.320 182.055 111.630 182.225 ;
        RECT 112.230 182.125 112.560 182.225 ;
        RECT 111.410 181.925 111.630 182.055 ;
        RECT 109.065 181.425 109.830 181.625 ;
        RECT 110.470 181.245 110.800 181.625 ;
        RECT 111.070 181.585 111.240 181.875 ;
        RECT 111.410 181.755 111.740 181.925 ;
        RECT 112.150 181.895 112.560 182.125 ;
        RECT 111.910 181.585 112.240 181.705 ;
        RECT 111.070 181.415 112.240 181.585 ;
        RECT 112.410 181.245 112.580 181.685 ;
        RECT 112.750 181.625 112.920 182.355 ;
        RECT 113.090 181.805 113.420 182.175 ;
        RECT 113.600 181.865 113.820 182.735 ;
        RECT 113.990 182.165 114.400 182.785 ;
        RECT 114.570 181.985 114.740 182.955 ;
        RECT 114.025 181.795 114.740 181.985 ;
        RECT 112.750 181.425 113.745 181.625 ;
        RECT 114.025 181.465 114.195 181.795 ;
        RECT 114.365 181.245 114.715 181.625 ;
        RECT 114.910 181.505 115.135 183.625 ;
        RECT 115.305 183.295 115.635 183.795 ;
        RECT 115.805 183.125 116.065 183.625 ;
        RECT 115.310 182.955 116.065 183.125 ;
        RECT 115.310 181.965 115.540 182.955 ;
        RECT 115.710 182.135 116.065 182.785 ;
        RECT 116.235 182.705 118.825 183.795 ;
        RECT 116.235 182.015 117.445 182.535 ;
        RECT 117.615 182.185 118.825 182.705 ;
        RECT 118.995 182.705 120.205 183.795 ;
        RECT 118.995 182.165 119.515 182.705 ;
        RECT 115.310 181.795 116.065 181.965 ;
        RECT 115.305 181.245 115.635 181.625 ;
        RECT 115.805 181.505 116.065 181.795 ;
        RECT 116.235 181.245 118.825 182.015 ;
        RECT 119.685 181.995 120.205 182.535 ;
        RECT 118.995 181.245 120.205 181.995 ;
        RECT 90.850 181.075 120.290 181.245 ;
        RECT 90.935 180.325 92.145 181.075 ;
        RECT 90.935 179.785 91.455 180.325 ;
        RECT 92.315 180.305 95.825 181.075 ;
        RECT 96.915 180.335 97.175 180.905 ;
        RECT 97.345 180.615 97.640 181.075 ;
        RECT 91.625 179.615 92.145 180.155 ;
        RECT 92.315 179.785 93.965 180.305 ;
        RECT 94.135 179.615 95.825 180.135 ;
        RECT 90.935 178.525 92.145 179.615 ;
        RECT 92.315 178.525 95.825 179.615 ;
        RECT 96.915 179.715 97.130 180.335 ;
        RECT 97.820 180.165 98.135 180.905 ;
        RECT 97.300 179.835 98.135 180.165 ;
        RECT 96.915 178.695 97.175 179.715 ;
        RECT 97.345 178.525 97.640 179.395 ;
        RECT 97.820 178.745 98.135 179.835 ;
        RECT 98.305 180.445 98.590 180.905 ;
        RECT 98.305 179.530 98.510 180.445 ;
        RECT 98.760 180.355 99.090 181.075 ;
        RECT 99.315 180.405 99.550 180.895 ;
        RECT 99.835 180.735 101.005 180.905 ;
        RECT 99.835 180.575 100.005 180.735 ;
        RECT 100.675 180.615 101.005 180.735 ;
        RECT 101.265 180.635 101.525 181.075 ;
        RECT 101.705 180.695 102.470 180.895 ;
        RECT 103.110 180.695 103.440 181.075 ;
        RECT 103.710 180.735 104.880 180.905 ;
        RECT 99.315 180.235 100.005 180.405 ;
        RECT 98.680 179.835 98.930 180.165 ;
        RECT 99.100 179.835 99.475 180.065 ;
        RECT 98.305 178.695 98.590 179.530 ;
        RECT 98.760 179.245 98.930 179.835 ;
        RECT 99.730 179.585 100.005 180.235 ;
        RECT 99.245 179.415 100.005 179.585 ;
        RECT 100.175 180.380 100.505 180.565 ;
        RECT 100.175 179.245 100.355 180.380 ;
        RECT 100.955 180.095 101.330 180.425 ;
        RECT 100.525 179.925 100.745 180.085 ;
        RECT 101.705 179.925 101.875 180.695 ;
        RECT 102.380 180.035 102.665 180.455 ;
        RECT 103.710 180.445 103.880 180.735 ;
        RECT 104.550 180.615 104.880 180.735 ;
        RECT 105.050 180.635 105.220 181.075 ;
        RECT 105.390 180.695 106.385 180.895 ;
        RECT 104.050 180.395 104.380 180.565 ;
        RECT 104.050 180.265 104.270 180.395 ;
        RECT 100.525 179.755 101.875 179.925 ;
        RECT 101.285 179.245 101.535 179.585 ;
        RECT 98.760 179.075 101.535 179.245 ;
        RECT 98.760 178.525 100.145 178.905 ;
        RECT 100.675 178.785 100.845 179.075 ;
        RECT 101.705 178.910 101.875 179.755 ;
        RECT 102.045 179.855 102.665 180.035 ;
        RECT 102.960 180.095 104.270 180.265 ;
        RECT 104.790 180.195 105.200 180.425 ;
        RECT 104.870 180.095 105.200 180.195 ;
        RECT 102.960 179.925 103.290 180.095 ;
        RECT 102.045 179.255 102.250 179.855 ;
        RECT 103.600 179.745 103.930 179.925 ;
        RECT 102.490 179.175 102.725 179.585 ;
        RECT 102.925 179.505 103.930 179.745 ;
        RECT 104.100 179.375 104.270 180.095 ;
        RECT 104.440 179.925 104.660 180.005 ;
        RECT 105.390 179.965 105.560 180.695 ;
        RECT 106.665 180.525 106.835 180.855 ;
        RECT 107.005 180.695 107.355 181.075 ;
        RECT 105.730 180.145 106.060 180.515 ;
        RECT 105.390 179.925 105.790 179.965 ;
        RECT 104.440 179.755 105.790 179.925 ;
        RECT 104.440 179.675 104.690 179.755 ;
        RECT 105.200 179.375 105.450 179.585 ;
        RECT 101.085 178.525 101.465 178.905 ;
        RECT 101.705 178.740 102.535 178.910 ;
        RECT 103.580 178.525 103.910 179.245 ;
        RECT 104.100 179.125 105.450 179.375 ;
        RECT 104.530 178.785 104.700 179.125 ;
        RECT 105.000 178.525 105.380 178.955 ;
        RECT 105.620 178.910 105.790 179.755 ;
        RECT 106.240 179.585 106.460 180.455 ;
        RECT 106.665 180.335 107.380 180.525 ;
        RECT 105.960 179.205 106.460 179.585 ;
        RECT 106.630 179.535 107.040 180.155 ;
        RECT 107.210 179.365 107.380 180.335 ;
        RECT 106.665 179.195 107.380 179.365 ;
        RECT 105.620 178.740 106.450 178.910 ;
        RECT 106.665 178.695 106.835 179.195 ;
        RECT 107.005 178.525 107.355 179.025 ;
        RECT 107.550 178.695 107.775 180.815 ;
        RECT 107.945 180.695 108.275 181.075 ;
        RECT 108.445 180.525 108.705 180.815 ;
        RECT 108.875 180.530 114.220 181.075 ;
        RECT 107.950 180.355 108.705 180.525 ;
        RECT 107.950 179.365 108.180 180.355 ;
        RECT 108.350 179.535 108.705 180.185 ;
        RECT 110.460 179.700 110.800 180.530 ;
        RECT 114.395 180.305 116.065 181.075 ;
        RECT 116.695 180.350 116.985 181.075 ;
        RECT 117.155 180.305 118.825 181.075 ;
        RECT 118.995 180.325 120.205 181.075 ;
        RECT 107.950 179.195 108.705 179.365 ;
        RECT 107.945 178.525 108.275 179.025 ;
        RECT 108.445 178.695 108.705 179.195 ;
        RECT 112.280 178.960 112.630 180.210 ;
        RECT 114.395 179.785 115.145 180.305 ;
        RECT 115.315 179.615 116.065 180.135 ;
        RECT 117.155 179.785 117.905 180.305 ;
        RECT 108.875 178.525 114.220 178.960 ;
        RECT 114.395 178.525 116.065 179.615 ;
        RECT 116.695 178.525 116.985 179.690 ;
        RECT 118.075 179.615 118.825 180.135 ;
        RECT 117.155 178.525 118.825 179.615 ;
        RECT 118.995 179.615 119.515 180.155 ;
        RECT 119.685 179.785 120.205 180.325 ;
        RECT 118.995 178.525 120.205 179.615 ;
        RECT 90.850 178.355 120.290 178.525 ;
        RECT 90.935 177.265 92.145 178.355 ;
        RECT 93.240 177.685 93.495 178.185 ;
        RECT 93.665 177.855 93.995 178.355 ;
        RECT 93.240 177.515 93.990 177.685 ;
        RECT 90.935 176.555 91.455 177.095 ;
        RECT 91.625 176.725 92.145 177.265 ;
        RECT 93.240 176.695 93.590 177.345 ;
        RECT 90.935 175.805 92.145 176.555 ;
        RECT 93.760 176.525 93.990 177.515 ;
        RECT 93.240 176.355 93.990 176.525 ;
        RECT 93.240 176.065 93.495 176.355 ;
        RECT 93.665 175.805 93.995 176.185 ;
        RECT 94.165 176.065 94.335 178.185 ;
        RECT 94.505 177.385 94.830 178.170 ;
        RECT 95.000 177.895 95.250 178.355 ;
        RECT 95.420 177.855 95.670 178.185 ;
        RECT 95.885 177.855 96.565 178.185 ;
        RECT 95.420 177.725 95.590 177.855 ;
        RECT 95.195 177.555 95.590 177.725 ;
        RECT 94.565 176.335 95.025 177.385 ;
        RECT 95.195 176.195 95.365 177.555 ;
        RECT 95.760 177.295 96.225 177.685 ;
        RECT 95.535 176.485 95.885 177.105 ;
        RECT 96.055 176.705 96.225 177.295 ;
        RECT 96.395 177.075 96.565 177.855 ;
        RECT 96.735 177.755 96.905 178.095 ;
        RECT 97.140 177.925 97.470 178.355 ;
        RECT 97.640 177.755 97.810 178.095 ;
        RECT 98.105 177.895 98.475 178.355 ;
        RECT 96.735 177.585 97.810 177.755 ;
        RECT 98.645 177.725 98.815 178.185 ;
        RECT 99.050 177.845 99.920 178.185 ;
        RECT 100.090 177.895 100.340 178.355 ;
        RECT 98.255 177.555 98.815 177.725 ;
        RECT 98.255 177.415 98.425 177.555 ;
        RECT 96.925 177.245 98.425 177.415 ;
        RECT 99.120 177.385 99.580 177.675 ;
        RECT 96.395 176.905 98.085 177.075 ;
        RECT 96.055 176.485 96.410 176.705 ;
        RECT 96.580 176.195 96.750 176.905 ;
        RECT 96.955 176.485 97.745 176.735 ;
        RECT 97.915 176.725 98.085 176.905 ;
        RECT 98.255 176.555 98.425 177.245 ;
        RECT 94.695 175.805 95.025 176.165 ;
        RECT 95.195 176.025 95.690 176.195 ;
        RECT 95.895 176.025 96.750 176.195 ;
        RECT 97.625 175.805 97.955 176.265 ;
        RECT 98.165 176.165 98.425 176.555 ;
        RECT 98.615 177.375 99.580 177.385 ;
        RECT 99.750 177.465 99.920 177.845 ;
        RECT 100.510 177.805 100.680 178.095 ;
        RECT 100.860 177.975 101.580 178.355 ;
        RECT 100.510 177.635 101.310 177.805 ;
        RECT 98.615 177.215 99.290 177.375 ;
        RECT 99.750 177.295 100.970 177.465 ;
        RECT 98.615 176.425 98.825 177.215 ;
        RECT 99.750 177.205 99.920 177.295 ;
        RECT 98.995 176.425 99.345 177.045 ;
        RECT 99.515 177.035 99.920 177.205 ;
        RECT 99.515 176.255 99.685 177.035 ;
        RECT 99.855 176.585 100.075 176.865 ;
        RECT 100.255 176.755 100.795 177.125 ;
        RECT 101.140 177.045 101.310 177.635 ;
        RECT 101.750 177.175 102.155 178.185 ;
        RECT 101.140 177.015 101.585 177.045 ;
        RECT 99.855 176.415 100.385 176.585 ;
        RECT 98.165 175.995 98.515 176.165 ;
        RECT 98.735 175.975 99.685 176.255 ;
        RECT 99.855 175.805 100.045 176.245 ;
        RECT 100.215 176.185 100.385 176.415 ;
        RECT 100.555 176.355 100.795 176.755 ;
        RECT 100.965 176.715 101.585 177.015 ;
        RECT 100.965 176.540 101.290 176.715 ;
        RECT 100.965 176.185 101.285 176.540 ;
        RECT 100.215 176.015 101.285 176.185 ;
        RECT 101.485 175.805 101.655 176.490 ;
        RECT 101.825 175.995 102.155 177.175 ;
        RECT 102.345 177.045 102.675 178.145 ;
        RECT 102.910 177.215 103.080 178.355 ;
        RECT 103.330 177.165 103.585 178.045 ;
        RECT 103.815 177.190 104.105 178.355 ;
        RECT 104.645 178.015 104.905 178.185 ;
        RECT 104.645 177.845 104.965 178.015 ;
        RECT 102.345 176.715 103.205 177.045 ;
        RECT 102.345 176.065 102.595 176.715 ;
        RECT 103.375 176.515 103.585 177.165 ;
        RECT 104.645 177.165 104.905 177.845 ;
        RECT 105.155 177.545 105.325 178.355 ;
        RECT 104.645 176.545 104.860 177.165 ;
        RECT 105.550 177.045 105.880 178.185 ;
        RECT 105.030 176.715 105.880 177.045 ;
        RECT 102.910 175.805 103.080 176.400 ;
        RECT 103.330 175.985 103.585 176.515 ;
        RECT 103.815 175.805 104.105 176.530 ;
        RECT 104.645 175.975 104.905 176.545 ;
        RECT 105.155 175.805 105.325 176.305 ;
        RECT 105.550 175.975 105.880 176.715 ;
        RECT 106.070 175.975 106.400 178.185 ;
        RECT 106.570 177.200 106.750 178.355 ;
        RECT 107.090 177.485 107.260 178.095 ;
        RECT 107.430 177.665 107.760 178.355 ;
        RECT 107.990 177.805 108.230 178.095 ;
        RECT 108.430 177.975 108.840 178.355 ;
        RECT 109.010 177.885 109.660 178.135 ;
        RECT 110.110 177.975 110.440 178.355 ;
        RECT 109.010 177.805 109.180 177.885 ;
        RECT 110.610 177.805 110.780 178.095 ;
        RECT 110.960 177.975 111.340 178.355 ;
        RECT 111.580 177.970 112.410 178.140 ;
        RECT 107.990 177.635 109.180 177.805 ;
        RECT 106.940 177.465 107.260 177.485 ;
        RECT 106.940 177.295 108.840 177.465 ;
        RECT 106.570 175.805 106.750 176.625 ;
        RECT 106.940 176.400 107.130 177.295 ;
        RECT 109.010 177.125 109.180 177.635 ;
        RECT 109.370 177.375 109.870 177.685 ;
        RECT 107.300 176.955 109.180 177.125 ;
        RECT 107.300 176.895 107.630 176.955 ;
        RECT 107.780 176.725 108.110 176.785 ;
        RECT 107.450 176.455 108.110 176.725 ;
        RECT 106.940 176.070 107.260 176.400 ;
        RECT 107.440 175.805 108.100 176.285 ;
        RECT 108.280 176.195 108.450 176.955 ;
        RECT 109.350 176.785 109.530 177.195 ;
        RECT 108.620 176.615 108.950 176.735 ;
        RECT 109.700 176.615 109.870 177.375 ;
        RECT 108.620 176.445 109.870 176.615 ;
        RECT 110.060 177.555 111.410 177.805 ;
        RECT 110.060 176.785 110.230 177.555 ;
        RECT 111.160 177.295 111.410 177.555 ;
        RECT 110.400 177.125 110.650 177.285 ;
        RECT 111.580 177.125 111.750 177.970 ;
        RECT 112.645 177.685 112.815 178.185 ;
        RECT 112.985 177.855 113.315 178.355 ;
        RECT 111.920 177.295 112.420 177.675 ;
        RECT 112.645 177.515 113.340 177.685 ;
        RECT 110.400 176.955 111.750 177.125 ;
        RECT 111.330 176.915 111.750 176.955 ;
        RECT 110.060 176.445 110.460 176.785 ;
        RECT 110.750 176.455 111.160 176.785 ;
        RECT 108.280 176.025 109.130 176.195 ;
        RECT 109.690 175.805 110.030 176.265 ;
        RECT 110.210 176.015 110.460 176.445 ;
        RECT 110.750 175.805 111.160 176.245 ;
        RECT 111.330 176.185 111.500 176.915 ;
        RECT 111.670 176.365 112.020 176.735 ;
        RECT 112.200 176.425 112.420 177.295 ;
        RECT 112.590 176.725 113.000 177.345 ;
        RECT 113.170 176.545 113.340 177.515 ;
        RECT 112.645 176.355 113.340 176.545 ;
        RECT 111.330 175.985 112.345 176.185 ;
        RECT 112.645 176.025 112.815 176.355 ;
        RECT 112.985 175.805 113.315 176.185 ;
        RECT 113.530 176.065 113.755 178.185 ;
        RECT 113.925 177.855 114.255 178.355 ;
        RECT 114.425 177.685 114.595 178.185 ;
        RECT 113.930 177.515 114.595 177.685 ;
        RECT 113.930 176.525 114.160 177.515 ;
        RECT 114.330 176.695 114.680 177.345 ;
        RECT 114.855 177.265 118.365 178.355 ;
        RECT 114.855 176.575 116.505 177.095 ;
        RECT 116.675 176.745 118.365 177.265 ;
        RECT 118.995 177.265 120.205 178.355 ;
        RECT 118.995 176.725 119.515 177.265 ;
        RECT 113.930 176.355 114.595 176.525 ;
        RECT 113.925 175.805 114.255 176.185 ;
        RECT 114.425 176.065 114.595 176.355 ;
        RECT 114.855 175.805 118.365 176.575 ;
        RECT 119.685 176.555 120.205 177.095 ;
        RECT 118.995 175.805 120.205 176.555 ;
        RECT 90.850 175.635 120.290 175.805 ;
        RECT 90.935 174.885 92.145 175.635 ;
        RECT 92.315 174.960 92.575 175.465 ;
        RECT 92.755 175.255 93.085 175.635 ;
        RECT 93.265 175.085 93.435 175.465 ;
        RECT 90.935 174.345 91.455 174.885 ;
        RECT 91.625 174.175 92.145 174.715 ;
        RECT 90.935 173.085 92.145 174.175 ;
        RECT 92.315 174.160 92.495 174.960 ;
        RECT 92.770 174.915 93.435 175.085 ;
        RECT 93.695 174.960 93.955 175.465 ;
        RECT 94.135 175.255 94.465 175.635 ;
        RECT 94.645 175.085 94.815 175.465 ;
        RECT 92.770 174.660 92.940 174.915 ;
        RECT 92.665 174.330 92.940 174.660 ;
        RECT 93.165 174.365 93.505 174.735 ;
        RECT 92.770 174.185 92.940 174.330 ;
        RECT 92.315 173.255 92.585 174.160 ;
        RECT 92.770 174.015 93.445 174.185 ;
        RECT 92.755 173.085 93.085 173.845 ;
        RECT 93.265 173.255 93.445 174.015 ;
        RECT 93.695 174.160 93.875 174.960 ;
        RECT 94.150 174.915 94.815 175.085 ;
        RECT 94.150 174.660 94.320 174.915 ;
        RECT 95.995 174.895 96.255 175.465 ;
        RECT 96.425 175.175 96.720 175.635 ;
        RECT 94.045 174.330 94.320 174.660 ;
        RECT 94.545 174.365 94.885 174.735 ;
        RECT 94.150 174.185 94.320 174.330 ;
        RECT 95.995 174.275 96.210 174.895 ;
        RECT 96.900 174.725 97.215 175.465 ;
        RECT 96.380 174.395 97.215 174.725 ;
        RECT 93.695 173.255 93.965 174.160 ;
        RECT 94.150 174.015 94.825 174.185 ;
        RECT 94.135 173.085 94.465 173.845 ;
        RECT 94.645 173.255 94.825 174.015 ;
        RECT 95.995 173.255 96.255 174.275 ;
        RECT 96.425 173.085 96.720 173.955 ;
        RECT 96.900 173.305 97.215 174.395 ;
        RECT 97.385 175.005 97.670 175.465 ;
        RECT 97.385 174.090 97.590 175.005 ;
        RECT 97.840 174.915 98.170 175.635 ;
        RECT 98.395 174.965 98.630 175.455 ;
        RECT 98.915 175.295 100.085 175.465 ;
        RECT 98.915 175.135 99.085 175.295 ;
        RECT 99.755 175.175 100.085 175.295 ;
        RECT 100.345 175.195 100.605 175.635 ;
        RECT 100.785 175.255 101.550 175.455 ;
        RECT 102.190 175.255 102.520 175.635 ;
        RECT 102.790 175.295 103.960 175.465 ;
        RECT 98.395 174.795 99.085 174.965 ;
        RECT 97.760 174.395 98.010 174.725 ;
        RECT 98.180 174.395 98.555 174.625 ;
        RECT 97.385 173.255 97.670 174.090 ;
        RECT 97.840 173.805 98.010 174.395 ;
        RECT 98.810 174.145 99.085 174.795 ;
        RECT 98.325 173.975 99.085 174.145 ;
        RECT 99.255 174.940 99.585 175.125 ;
        RECT 99.255 173.805 99.435 174.940 ;
        RECT 100.035 174.655 100.410 174.985 ;
        RECT 99.605 174.485 99.825 174.645 ;
        RECT 100.785 174.485 100.955 175.255 ;
        RECT 101.460 174.595 101.745 175.015 ;
        RECT 102.790 175.005 102.960 175.295 ;
        RECT 103.630 175.175 103.960 175.295 ;
        RECT 104.130 175.195 104.300 175.635 ;
        RECT 104.470 175.255 105.465 175.455 ;
        RECT 103.130 174.955 103.460 175.125 ;
        RECT 103.130 174.825 103.350 174.955 ;
        RECT 99.605 174.315 100.955 174.485 ;
        RECT 100.365 173.805 100.615 174.145 ;
        RECT 97.840 173.635 100.615 173.805 ;
        RECT 97.840 173.085 99.225 173.465 ;
        RECT 99.755 173.345 99.925 173.635 ;
        RECT 100.785 173.470 100.955 174.315 ;
        RECT 101.125 174.415 101.745 174.595 ;
        RECT 102.040 174.655 103.350 174.825 ;
        RECT 103.870 174.755 104.280 174.985 ;
        RECT 103.950 174.655 104.280 174.755 ;
        RECT 102.040 174.485 102.370 174.655 ;
        RECT 101.125 173.815 101.330 174.415 ;
        RECT 102.680 174.305 103.010 174.485 ;
        RECT 101.570 173.735 101.805 174.145 ;
        RECT 102.005 174.065 103.010 174.305 ;
        RECT 103.180 173.935 103.350 174.655 ;
        RECT 103.520 174.485 103.740 174.565 ;
        RECT 104.470 174.525 104.640 175.255 ;
        RECT 105.745 175.085 105.915 175.415 ;
        RECT 106.085 175.255 106.435 175.635 ;
        RECT 104.810 174.705 105.140 175.075 ;
        RECT 104.470 174.485 104.870 174.525 ;
        RECT 103.520 174.315 104.870 174.485 ;
        RECT 103.520 174.235 103.770 174.315 ;
        RECT 104.280 173.935 104.530 174.145 ;
        RECT 100.165 173.085 100.545 173.465 ;
        RECT 100.785 173.300 101.615 173.470 ;
        RECT 102.660 173.085 102.990 173.805 ;
        RECT 103.180 173.685 104.530 173.935 ;
        RECT 103.610 173.345 103.780 173.685 ;
        RECT 104.080 173.085 104.460 173.515 ;
        RECT 104.700 173.470 104.870 174.315 ;
        RECT 105.320 174.145 105.540 175.015 ;
        RECT 105.745 174.895 106.460 175.085 ;
        RECT 105.040 173.765 105.540 174.145 ;
        RECT 105.710 174.095 106.120 174.715 ;
        RECT 106.290 173.925 106.460 174.895 ;
        RECT 105.745 173.755 106.460 173.925 ;
        RECT 104.700 173.300 105.530 173.470 ;
        RECT 105.745 173.255 105.915 173.755 ;
        RECT 106.085 173.085 106.435 173.585 ;
        RECT 106.630 173.255 106.855 175.375 ;
        RECT 107.025 175.255 107.355 175.635 ;
        RECT 107.525 175.085 107.785 175.375 ;
        RECT 107.955 175.090 113.300 175.635 ;
        RECT 107.030 174.915 107.785 175.085 ;
        RECT 107.030 173.925 107.260 174.915 ;
        RECT 107.430 174.095 107.785 174.745 ;
        RECT 109.540 174.260 109.880 175.090 ;
        RECT 113.475 174.865 116.065 175.635 ;
        RECT 116.695 174.910 116.985 175.635 ;
        RECT 117.155 174.865 118.825 175.635 ;
        RECT 118.995 174.885 120.205 175.635 ;
        RECT 107.030 173.755 107.785 173.925 ;
        RECT 107.025 173.085 107.355 173.585 ;
        RECT 107.525 173.255 107.785 173.755 ;
        RECT 111.360 173.520 111.710 174.770 ;
        RECT 113.475 174.345 114.685 174.865 ;
        RECT 114.855 174.175 116.065 174.695 ;
        RECT 117.155 174.345 117.905 174.865 ;
        RECT 107.955 173.085 113.300 173.520 ;
        RECT 113.475 173.085 116.065 174.175 ;
        RECT 116.695 173.085 116.985 174.250 ;
        RECT 118.075 174.175 118.825 174.695 ;
        RECT 117.155 173.085 118.825 174.175 ;
        RECT 118.995 174.175 119.515 174.715 ;
        RECT 119.685 174.345 120.205 174.885 ;
        RECT 118.995 173.085 120.205 174.175 ;
        RECT 90.850 172.915 120.290 173.085 ;
        RECT 90.935 171.825 92.145 172.915 ;
        RECT 92.405 172.170 92.675 172.915 ;
        RECT 93.305 172.910 99.580 172.915 ;
        RECT 92.845 172.000 93.135 172.740 ;
        RECT 93.305 172.185 93.560 172.910 ;
        RECT 93.745 172.015 94.005 172.740 ;
        RECT 94.175 172.185 94.420 172.910 ;
        RECT 94.605 172.015 94.865 172.740 ;
        RECT 95.035 172.185 95.280 172.910 ;
        RECT 95.465 172.015 95.725 172.740 ;
        RECT 95.895 172.185 96.140 172.910 ;
        RECT 96.310 172.015 96.570 172.740 ;
        RECT 96.740 172.185 97.000 172.910 ;
        RECT 97.170 172.015 97.430 172.740 ;
        RECT 97.600 172.185 97.860 172.910 ;
        RECT 98.030 172.015 98.290 172.740 ;
        RECT 98.460 172.185 98.720 172.910 ;
        RECT 98.890 172.015 99.150 172.740 ;
        RECT 99.320 172.115 99.580 172.910 ;
        RECT 93.745 172.000 99.150 172.015 ;
        RECT 90.935 171.115 91.455 171.655 ;
        RECT 91.625 171.285 92.145 171.825 ;
        RECT 92.405 171.775 99.150 172.000 ;
        RECT 92.405 171.185 93.570 171.775 ;
        RECT 99.750 171.605 100.000 172.740 ;
        RECT 100.180 172.105 100.440 172.915 ;
        RECT 100.615 171.605 100.860 172.745 ;
        RECT 101.040 172.105 101.335 172.915 ;
        RECT 102.435 171.840 102.705 172.745 ;
        RECT 102.875 172.155 103.205 172.915 ;
        RECT 103.385 171.985 103.565 172.745 ;
        RECT 93.740 171.355 100.860 171.605 ;
        RECT 90.935 170.365 92.145 171.115 ;
        RECT 92.405 171.015 99.150 171.185 ;
        RECT 92.405 170.365 92.705 170.845 ;
        RECT 92.875 170.560 93.135 171.015 ;
        RECT 93.305 170.365 93.565 170.845 ;
        RECT 93.745 170.560 94.005 171.015 ;
        RECT 94.175 170.365 94.425 170.845 ;
        RECT 94.605 170.560 94.865 171.015 ;
        RECT 95.035 170.365 95.285 170.845 ;
        RECT 95.465 170.560 95.725 171.015 ;
        RECT 95.895 170.365 96.140 170.845 ;
        RECT 96.310 170.560 96.585 171.015 ;
        RECT 96.755 170.365 97.000 170.845 ;
        RECT 97.170 170.560 97.430 171.015 ;
        RECT 97.600 170.365 97.860 170.845 ;
        RECT 98.030 170.560 98.290 171.015 ;
        RECT 98.460 170.365 98.720 170.845 ;
        RECT 98.890 170.560 99.150 171.015 ;
        RECT 99.320 170.365 99.580 170.925 ;
        RECT 99.750 170.545 100.000 171.355 ;
        RECT 100.180 170.365 100.440 170.890 ;
        RECT 100.610 170.545 100.860 171.355 ;
        RECT 101.030 171.045 101.345 171.605 ;
        RECT 102.435 171.040 102.615 171.840 ;
        RECT 102.890 171.815 103.565 171.985 ;
        RECT 102.890 171.670 103.060 171.815 ;
        RECT 103.815 171.750 104.105 172.915 ;
        RECT 104.365 172.170 104.635 172.915 ;
        RECT 105.265 172.910 111.540 172.915 ;
        RECT 104.805 172.000 105.095 172.740 ;
        RECT 105.265 172.185 105.520 172.910 ;
        RECT 105.705 172.015 105.965 172.740 ;
        RECT 106.135 172.185 106.380 172.910 ;
        RECT 106.565 172.015 106.825 172.740 ;
        RECT 106.995 172.185 107.240 172.910 ;
        RECT 107.425 172.015 107.685 172.740 ;
        RECT 107.855 172.185 108.100 172.910 ;
        RECT 108.270 172.015 108.530 172.740 ;
        RECT 108.700 172.185 108.960 172.910 ;
        RECT 109.130 172.015 109.390 172.740 ;
        RECT 109.560 172.185 109.820 172.910 ;
        RECT 109.990 172.015 110.250 172.740 ;
        RECT 110.420 172.185 110.680 172.910 ;
        RECT 110.850 172.015 111.110 172.740 ;
        RECT 111.280 172.115 111.540 172.910 ;
        RECT 105.705 172.000 111.110 172.015 ;
        RECT 104.365 171.775 111.110 172.000 ;
        RECT 102.785 171.340 103.060 171.670 ;
        RECT 102.890 171.085 103.060 171.340 ;
        RECT 103.285 171.265 103.625 171.635 ;
        RECT 104.365 171.185 105.530 171.775 ;
        RECT 111.710 171.605 111.960 172.740 ;
        RECT 112.140 172.105 112.400 172.915 ;
        RECT 112.575 171.605 112.820 172.745 ;
        RECT 113.000 172.105 113.295 172.915 ;
        RECT 113.475 171.825 116.065 172.915 ;
        RECT 105.700 171.355 112.820 171.605 ;
        RECT 101.040 170.365 101.345 170.875 ;
        RECT 102.435 170.535 102.695 171.040 ;
        RECT 102.890 170.915 103.555 171.085 ;
        RECT 102.875 170.365 103.205 170.745 ;
        RECT 103.385 170.535 103.555 170.915 ;
        RECT 103.815 170.365 104.105 171.090 ;
        RECT 104.365 171.015 111.110 171.185 ;
        RECT 104.365 170.365 104.665 170.845 ;
        RECT 104.835 170.560 105.095 171.015 ;
        RECT 105.265 170.365 105.525 170.845 ;
        RECT 105.705 170.560 105.965 171.015 ;
        RECT 106.135 170.365 106.385 170.845 ;
        RECT 106.565 170.560 106.825 171.015 ;
        RECT 106.995 170.365 107.245 170.845 ;
        RECT 107.425 170.560 107.685 171.015 ;
        RECT 107.855 170.365 108.100 170.845 ;
        RECT 108.270 170.560 108.545 171.015 ;
        RECT 108.715 170.365 108.960 170.845 ;
        RECT 109.130 170.560 109.390 171.015 ;
        RECT 109.560 170.365 109.820 170.845 ;
        RECT 109.990 170.560 110.250 171.015 ;
        RECT 110.420 170.365 110.680 170.845 ;
        RECT 110.850 170.560 111.110 171.015 ;
        RECT 111.280 170.365 111.540 170.925 ;
        RECT 111.710 170.545 111.960 171.355 ;
        RECT 112.140 170.365 112.400 170.890 ;
        RECT 112.570 170.545 112.820 171.355 ;
        RECT 112.990 171.045 113.305 171.605 ;
        RECT 113.475 171.135 114.685 171.655 ;
        RECT 114.855 171.305 116.065 171.825 ;
        RECT 116.695 171.750 116.985 172.915 ;
        RECT 117.155 171.825 118.825 172.915 ;
        RECT 117.155 171.135 117.905 171.655 ;
        RECT 118.075 171.305 118.825 171.825 ;
        RECT 118.995 171.825 120.205 172.915 ;
        RECT 118.995 171.285 119.515 171.825 ;
        RECT 113.000 170.365 113.305 170.875 ;
        RECT 113.475 170.365 116.065 171.135 ;
        RECT 116.695 170.365 116.985 171.090 ;
        RECT 117.155 170.365 118.825 171.135 ;
        RECT 119.685 171.115 120.205 171.655 ;
        RECT 118.995 170.365 120.205 171.115 ;
        RECT 90.850 170.195 120.290 170.365 ;
        RECT 47.465 153.445 48.665 153.450 ;
        RECT 47.465 152.835 52.595 153.445 ;
        RECT 54.080 152.840 59.300 153.445 ;
        RECT 47.465 150.585 49.025 152.835 ;
        RECT 49.695 152.275 51.735 152.445 ;
        RECT 49.355 151.215 49.525 152.215 ;
        RECT 51.905 151.215 52.075 152.215 ;
        RECT 49.695 150.985 51.735 151.155 ;
        RECT 52.415 150.585 52.585 152.835 ;
        RECT 47.465 150.415 52.585 150.585 ;
        RECT 47.465 147.085 49.025 150.415 ;
        RECT 49.695 149.845 51.735 150.015 ;
        RECT 49.355 149.285 49.525 149.785 ;
        RECT 51.905 149.285 52.075 149.785 ;
        RECT 49.695 149.055 51.735 149.225 ;
        RECT 49.355 148.495 49.525 148.995 ;
        RECT 51.905 148.495 52.075 148.995 ;
        RECT 49.695 148.265 51.735 148.435 ;
        RECT 49.355 147.705 49.525 148.205 ;
        RECT 51.905 147.705 52.075 148.205 ;
        RECT 49.695 147.475 51.735 147.645 ;
        RECT 52.415 147.085 52.585 150.415 ;
        RECT 54.085 150.585 54.255 152.840 ;
        RECT 54.980 152.275 57.020 152.445 ;
        RECT 54.595 151.215 54.765 152.215 ;
        RECT 57.235 151.215 57.405 152.215 ;
        RECT 54.980 150.985 57.020 151.155 ;
        RECT 57.740 150.585 59.300 152.840 ;
        RECT 54.085 150.415 59.300 150.585 ;
        RECT 47.465 146.630 52.590 147.085 ;
        RECT 54.085 145.500 54.255 150.415 ;
        RECT 54.980 149.845 57.020 150.015 ;
        RECT 54.595 149.285 54.765 149.785 ;
        RECT 57.235 149.285 57.405 149.785 ;
        RECT 54.980 149.055 57.020 149.225 ;
        RECT 54.595 148.495 54.765 148.995 ;
        RECT 57.235 148.495 57.405 148.995 ;
        RECT 54.980 148.265 57.020 148.435 ;
        RECT 54.595 147.705 54.765 148.205 ;
        RECT 57.235 147.705 57.405 148.205 ;
        RECT 54.980 147.475 57.020 147.645 ;
        RECT 54.595 146.915 54.765 147.415 ;
        RECT 57.235 146.915 57.405 147.415 ;
        RECT 54.980 146.685 57.020 146.855 ;
        RECT 54.595 146.125 54.765 146.625 ;
        RECT 57.235 146.125 57.405 146.625 ;
        RECT 54.980 145.895 57.020 146.065 ;
        RECT 57.740 145.500 59.300 150.415 ;
        RECT 60.995 153.420 62.195 153.425 ;
        RECT 74.800 153.420 76.000 153.425 ;
        RECT 88.490 153.420 89.690 153.425 ;
        RECT 60.995 152.810 66.125 153.420 ;
        RECT 67.610 152.815 72.830 153.420 ;
        RECT 60.995 150.560 62.555 152.810 ;
        RECT 63.225 152.250 65.265 152.420 ;
        RECT 62.885 151.190 63.055 152.190 ;
        RECT 65.435 151.190 65.605 152.190 ;
        RECT 63.225 150.960 65.265 151.130 ;
        RECT 65.945 150.560 66.115 152.810 ;
        RECT 60.995 150.390 66.115 150.560 ;
        RECT 60.995 147.060 62.555 150.390 ;
        RECT 63.225 149.820 65.265 149.990 ;
        RECT 62.885 149.260 63.055 149.760 ;
        RECT 65.435 149.260 65.605 149.760 ;
        RECT 63.225 149.030 65.265 149.200 ;
        RECT 62.885 148.470 63.055 148.970 ;
        RECT 65.435 148.470 65.605 148.970 ;
        RECT 63.225 148.240 65.265 148.410 ;
        RECT 62.885 147.680 63.055 148.180 ;
        RECT 65.435 147.680 65.605 148.180 ;
        RECT 63.225 147.450 65.265 147.620 ;
        RECT 65.945 147.060 66.115 150.390 ;
        RECT 67.615 150.560 67.785 152.815 ;
        RECT 68.510 152.250 70.550 152.420 ;
        RECT 68.125 151.190 68.295 152.190 ;
        RECT 70.765 151.190 70.935 152.190 ;
        RECT 68.510 150.960 70.550 151.130 ;
        RECT 71.270 150.560 72.830 152.815 ;
        RECT 67.615 150.390 72.830 150.560 ;
        RECT 60.995 146.605 66.120 147.060 ;
        RECT 54.080 144.955 59.300 145.500 ;
        RECT 67.615 145.475 67.785 150.390 ;
        RECT 68.510 149.820 70.550 149.990 ;
        RECT 68.125 149.260 68.295 149.760 ;
        RECT 70.765 149.260 70.935 149.760 ;
        RECT 68.510 149.030 70.550 149.200 ;
        RECT 68.125 148.470 68.295 148.970 ;
        RECT 70.765 148.470 70.935 148.970 ;
        RECT 68.510 148.240 70.550 148.410 ;
        RECT 68.125 147.680 68.295 148.180 ;
        RECT 70.765 147.680 70.935 148.180 ;
        RECT 68.510 147.450 70.550 147.620 ;
        RECT 68.125 146.890 68.295 147.390 ;
        RECT 70.765 146.890 70.935 147.390 ;
        RECT 68.510 146.660 70.550 146.830 ;
        RECT 68.125 146.100 68.295 146.600 ;
        RECT 70.765 146.100 70.935 146.600 ;
        RECT 68.510 145.870 70.550 146.040 ;
        RECT 71.270 145.475 72.830 150.390 ;
        RECT 74.800 152.810 79.930 153.420 ;
        RECT 81.415 152.815 86.635 153.420 ;
        RECT 74.800 150.560 76.360 152.810 ;
        RECT 77.030 152.250 79.070 152.420 ;
        RECT 76.690 151.190 76.860 152.190 ;
        RECT 79.240 151.190 79.410 152.190 ;
        RECT 77.030 150.960 79.070 151.130 ;
        RECT 79.750 150.560 79.920 152.810 ;
        RECT 74.800 150.390 79.920 150.560 ;
        RECT 74.800 147.060 76.360 150.390 ;
        RECT 77.030 149.820 79.070 149.990 ;
        RECT 76.690 149.260 76.860 149.760 ;
        RECT 79.240 149.260 79.410 149.760 ;
        RECT 77.030 149.030 79.070 149.200 ;
        RECT 76.690 148.470 76.860 148.970 ;
        RECT 79.240 148.470 79.410 148.970 ;
        RECT 77.030 148.240 79.070 148.410 ;
        RECT 76.690 147.680 76.860 148.180 ;
        RECT 79.240 147.680 79.410 148.180 ;
        RECT 77.030 147.450 79.070 147.620 ;
        RECT 79.750 147.060 79.920 150.390 ;
        RECT 81.420 150.560 81.590 152.815 ;
        RECT 82.315 152.250 84.355 152.420 ;
        RECT 81.930 151.190 82.100 152.190 ;
        RECT 84.570 151.190 84.740 152.190 ;
        RECT 82.315 150.960 84.355 151.130 ;
        RECT 85.075 150.560 86.635 152.815 ;
        RECT 81.420 150.390 86.635 150.560 ;
        RECT 74.800 146.605 79.925 147.060 ;
        RECT 81.420 145.475 81.590 150.390 ;
        RECT 82.315 149.820 84.355 149.990 ;
        RECT 81.930 149.260 82.100 149.760 ;
        RECT 84.570 149.260 84.740 149.760 ;
        RECT 82.315 149.030 84.355 149.200 ;
        RECT 81.930 148.470 82.100 148.970 ;
        RECT 84.570 148.470 84.740 148.970 ;
        RECT 82.315 148.240 84.355 148.410 ;
        RECT 81.930 147.680 82.100 148.180 ;
        RECT 84.570 147.680 84.740 148.180 ;
        RECT 82.315 147.450 84.355 147.620 ;
        RECT 81.930 146.890 82.100 147.390 ;
        RECT 84.570 146.890 84.740 147.390 ;
        RECT 82.315 146.660 84.355 146.830 ;
        RECT 81.930 146.100 82.100 146.600 ;
        RECT 84.570 146.100 84.740 146.600 ;
        RECT 82.315 145.870 84.355 146.040 ;
        RECT 85.075 145.475 86.635 150.390 ;
        RECT 88.490 152.810 93.620 153.420 ;
        RECT 95.105 152.815 100.325 153.420 ;
        RECT 88.490 150.560 90.050 152.810 ;
        RECT 90.720 152.250 92.760 152.420 ;
        RECT 90.380 151.190 90.550 152.190 ;
        RECT 92.930 151.190 93.100 152.190 ;
        RECT 90.720 150.960 92.760 151.130 ;
        RECT 93.440 150.560 93.610 152.810 ;
        RECT 88.490 150.390 93.610 150.560 ;
        RECT 88.490 147.060 90.050 150.390 ;
        RECT 90.720 149.820 92.760 149.990 ;
        RECT 90.380 149.260 90.550 149.760 ;
        RECT 92.930 149.260 93.100 149.760 ;
        RECT 90.720 149.030 92.760 149.200 ;
        RECT 90.380 148.470 90.550 148.970 ;
        RECT 92.930 148.470 93.100 148.970 ;
        RECT 90.720 148.240 92.760 148.410 ;
        RECT 90.380 147.680 90.550 148.180 ;
        RECT 92.930 147.680 93.100 148.180 ;
        RECT 90.720 147.450 92.760 147.620 ;
        RECT 93.440 147.060 93.610 150.390 ;
        RECT 95.110 150.560 95.280 152.815 ;
        RECT 96.005 152.250 98.045 152.420 ;
        RECT 95.620 151.190 95.790 152.190 ;
        RECT 98.260 151.190 98.430 152.190 ;
        RECT 96.005 150.960 98.045 151.130 ;
        RECT 98.765 150.560 100.325 152.815 ;
        RECT 95.110 150.390 100.325 150.560 ;
        RECT 88.490 146.605 93.615 147.060 ;
        RECT 95.110 145.475 95.280 150.390 ;
        RECT 96.005 149.820 98.045 149.990 ;
        RECT 95.620 149.260 95.790 149.760 ;
        RECT 98.260 149.260 98.430 149.760 ;
        RECT 96.005 149.030 98.045 149.200 ;
        RECT 95.620 148.470 95.790 148.970 ;
        RECT 98.260 148.470 98.430 148.970 ;
        RECT 96.005 148.240 98.045 148.410 ;
        RECT 95.620 147.680 95.790 148.180 ;
        RECT 98.260 147.680 98.430 148.180 ;
        RECT 96.005 147.450 98.045 147.620 ;
        RECT 95.620 146.890 95.790 147.390 ;
        RECT 98.260 146.890 98.430 147.390 ;
        RECT 96.005 146.660 98.045 146.830 ;
        RECT 95.620 146.100 95.790 146.600 ;
        RECT 98.260 146.100 98.430 146.600 ;
        RECT 96.005 145.870 98.045 146.040 ;
        RECT 98.765 145.475 100.325 150.390 ;
        RECT 67.610 144.930 72.830 145.475 ;
        RECT 81.415 144.930 86.635 145.475 ;
        RECT 95.105 144.930 100.325 145.475 ;
        RECT 66.585 138.565 68.235 138.735 ;
        RECT 66.585 138.265 66.755 138.565 ;
        RECT 66.200 138.015 66.765 138.265 ;
        RECT 67.235 138.015 67.585 138.085 ;
        RECT 66.200 135.990 67.585 138.015 ;
        RECT 68.065 136.945 68.235 138.565 ;
        RECT 66.200 121.455 66.765 135.990 ;
        RECT 67.235 135.925 67.585 135.990 ;
        RECT 68.050 136.935 68.770 136.945 ;
        RECT 68.050 136.765 70.240 136.935 ;
        RECT 67.235 121.925 67.585 124.085 ;
        RECT 68.050 121.455 68.770 136.765 ;
        RECT 70.070 136.545 70.240 136.765 ;
        RECT 76.090 136.735 76.525 136.740 ;
        RECT 74.620 136.565 76.525 136.735 ;
        RECT 70.050 136.535 70.780 136.545 ;
        RECT 72.070 136.535 72.790 136.545 ;
        RECT 74.620 136.540 74.790 136.565 ;
        RECT 74.085 136.535 74.790 136.540 ;
        RECT 70.050 136.395 74.790 136.535 ;
        RECT 70.050 136.365 74.800 136.395 ;
        RECT 69.240 134.125 69.590 136.285 ;
        RECT 69.240 121.925 69.590 124.085 ;
        RECT 70.050 121.455 70.780 136.365 ;
        RECT 71.250 133.725 71.600 135.885 ;
        RECT 71.250 121.925 71.600 124.085 ;
        RECT 72.070 121.455 72.790 136.365 ;
        RECT 73.260 133.725 73.610 135.885 ;
        RECT 73.260 121.925 73.610 124.085 ;
        RECT 74.085 121.455 74.800 136.365 ;
        RECT 75.270 133.925 75.620 136.085 ;
        RECT 75.270 121.925 75.620 124.085 ;
        RECT 76.090 121.455 76.525 136.565 ;
        RECT 85.315 136.325 114.315 137.700 ;
        RECT 85.320 130.945 87.485 136.325 ;
        RECT 88.065 135.835 92.065 136.005 ;
        RECT 87.835 131.625 88.005 135.665 ;
        RECT 92.125 131.625 92.295 135.665 ;
        RECT 88.065 131.285 92.065 131.455 ;
        RECT 92.695 130.945 92.865 136.325 ;
        RECT 93.495 135.835 97.495 136.005 ;
        RECT 93.265 131.625 93.435 135.665 ;
        RECT 97.555 131.625 97.725 135.665 ;
        RECT 93.495 131.285 97.495 131.455 ;
        RECT 98.105 131.110 100.390 136.325 ;
        RECT 101.025 135.800 103.065 135.970 ;
        RECT 100.685 131.740 100.855 135.740 ;
        RECT 103.235 131.740 103.405 135.740 ;
        RECT 101.025 131.510 103.065 131.680 ;
        RECT 103.745 131.110 103.915 136.325 ;
        RECT 104.595 135.800 106.635 135.970 ;
        RECT 104.255 131.740 104.425 135.740 ;
        RECT 106.805 131.740 106.975 135.740 ;
        RECT 107.290 134.235 114.310 136.325 ;
        RECT 107.290 132.390 110.285 134.235 ;
        RECT 110.885 133.850 111.385 134.020 ;
        RECT 110.655 133.030 110.825 133.680 ;
        RECT 111.445 133.030 111.615 133.680 ;
        RECT 110.885 132.690 111.385 132.860 ;
        RECT 111.995 132.390 114.310 134.235 ;
        RECT 104.595 131.510 106.635 131.680 ;
        RECT 107.290 131.110 114.325 132.390 ;
        RECT 98.105 130.945 114.325 131.110 ;
        RECT 85.320 130.940 114.325 130.945 ;
        RECT 85.320 130.775 100.390 130.940 ;
        RECT 85.320 130.570 87.485 130.775 ;
        RECT 98.105 130.590 100.390 130.775 ;
        RECT 107.290 130.630 114.325 130.940 ;
        RECT 107.290 130.610 110.285 130.630 ;
        RECT 85.845 128.195 87.015 128.200 ;
        RECT 66.200 121.430 76.525 121.455 ;
        RECT 85.300 128.010 87.440 128.195 ;
        RECT 94.100 128.010 96.505 128.195 ;
        RECT 85.300 128.005 96.505 128.010 ;
        RECT 107.730 128.190 110.245 128.195 ;
        RECT 107.730 128.005 114.310 128.190 ;
        RECT 85.300 127.840 114.310 128.005 ;
        RECT 85.300 122.360 87.440 127.840 ;
        RECT 88.070 127.330 90.070 127.500 ;
        RECT 87.840 123.075 88.010 127.115 ;
        RECT 90.130 123.075 90.300 127.115 ;
        RECT 88.070 122.690 90.070 122.860 ;
        RECT 90.700 122.360 90.870 127.840 ;
        RECT 94.100 127.835 114.310 127.840 ;
        RECT 91.500 127.330 93.500 127.500 ;
        RECT 91.270 123.075 91.440 127.115 ;
        RECT 93.560 123.075 93.730 127.115 ;
        RECT 91.500 122.690 93.500 122.860 ;
        RECT 94.100 122.360 96.505 127.835 ;
        RECT 97.115 127.325 99.115 127.495 ;
        RECT 99.405 127.325 101.405 127.495 ;
        RECT 96.885 123.070 97.055 127.110 ;
        RECT 99.175 123.070 99.345 127.110 ;
        RECT 101.465 123.070 101.635 127.110 ;
        RECT 97.115 122.685 99.115 122.855 ;
        RECT 99.405 122.685 101.405 122.855 ;
        RECT 102.035 122.360 102.205 127.835 ;
        RECT 102.835 127.325 104.835 127.495 ;
        RECT 105.125 127.325 107.125 127.495 ;
        RECT 102.605 123.070 102.775 127.110 ;
        RECT 104.895 123.070 105.065 127.110 ;
        RECT 107.185 123.070 107.355 127.110 ;
        RECT 107.730 126.790 114.310 127.835 ;
        RECT 107.730 124.860 110.245 126.790 ;
        RECT 110.860 126.320 111.360 126.490 ;
        RECT 110.630 125.565 110.800 126.105 ;
        RECT 111.420 125.565 111.590 126.105 ;
        RECT 110.860 125.180 111.360 125.350 ;
        RECT 111.975 124.860 114.310 126.790 ;
        RECT 102.835 122.685 104.835 122.855 ;
        RECT 105.125 122.685 107.125 122.855 ;
        RECT 107.725 122.360 114.310 124.860 ;
        RECT 119.290 124.620 125.370 125.085 ;
        RECT 66.200 121.045 76.520 121.430 ;
        RECT 66.200 120.735 74.680 121.045 ;
        RECT 85.300 120.860 114.315 122.360 ;
        RECT 112.250 120.850 114.315 120.860 ;
        RECT 66.200 110.830 68.770 120.735 ;
        RECT 69.240 118.105 69.590 120.265 ;
        RECT 69.240 111.305 69.590 113.465 ;
        RECT 70.060 110.830 70.780 120.735 ;
        RECT 71.250 118.105 71.600 120.265 ;
        RECT 71.250 111.305 71.600 113.465 ;
        RECT 72.070 110.830 72.790 120.735 ;
        RECT 73.260 118.105 73.610 120.265 ;
        RECT 73.260 111.305 73.610 113.465 ;
        RECT 74.085 110.830 74.680 120.735 ;
        RECT 119.290 119.140 119.715 124.620 ;
        RECT 120.335 124.120 121.335 124.290 ;
        RECT 120.105 119.865 120.275 123.905 ;
        RECT 121.395 119.865 121.565 123.905 ;
        RECT 121.955 121.610 125.370 124.620 ;
        RECT 120.335 119.480 121.335 119.650 ;
        RECT 121.955 119.140 122.675 121.610 ;
        RECT 123.295 121.120 124.295 121.290 ;
        RECT 123.065 119.865 123.235 120.905 ;
        RECT 124.355 119.865 124.525 120.905 ;
        RECT 123.295 119.480 124.295 119.650 ;
        RECT 124.915 119.140 125.370 121.610 ;
        RECT 119.290 118.970 125.370 119.140 ;
        RECT 119.290 118.955 119.715 118.970 ;
        RECT 121.955 118.955 122.675 118.970 ;
        RECT 124.915 118.955 125.370 118.970 ;
        RECT 119.285 117.300 119.710 117.305 ;
        RECT 121.950 117.300 122.670 117.305 ;
        RECT 124.900 117.300 125.370 117.305 ;
        RECT 119.285 117.130 125.370 117.300 ;
        RECT 66.200 110.765 74.680 110.830 ;
        RECT 81.750 114.135 106.100 115.810 ;
        RECT 66.200 110.200 74.675 110.765 ;
        RECT 81.750 108.660 82.585 114.135 ;
        RECT 83.200 113.640 85.200 113.810 ;
        RECT 82.970 109.385 83.140 113.425 ;
        RECT 85.260 113.350 85.430 113.425 ;
        RECT 85.825 113.350 89.530 114.135 ;
        RECT 90.150 113.640 91.150 113.810 ;
        RECT 85.255 111.405 89.530 113.350 ;
        RECT 85.260 109.385 85.430 111.405 ;
        RECT 83.200 109.000 85.200 109.170 ;
        RECT 85.830 108.660 86.000 111.405 ;
        RECT 81.750 108.490 86.000 108.660 ;
        RECT 89.350 108.660 89.520 111.405 ;
        RECT 89.920 109.385 90.090 113.425 ;
        RECT 91.210 109.385 91.380 113.425 ;
        RECT 90.150 109.000 91.150 109.170 ;
        RECT 91.780 108.660 91.950 114.135 ;
        RECT 92.580 113.640 93.580 113.810 ;
        RECT 92.350 109.385 92.520 113.425 ;
        RECT 93.640 109.385 93.810 113.425 ;
        RECT 94.200 113.355 97.920 114.135 ;
        RECT 98.540 113.645 100.540 113.815 ;
        RECT 98.310 113.355 98.480 113.430 ;
        RECT 94.200 111.405 98.490 113.355 ;
        RECT 92.580 109.000 93.580 109.170 ;
        RECT 94.210 108.660 94.380 111.405 ;
        RECT 89.350 108.490 94.380 108.660 ;
        RECT 97.740 108.665 97.910 111.405 ;
        RECT 98.310 109.390 98.480 111.405 ;
        RECT 100.600 109.390 100.770 113.430 ;
        RECT 101.160 111.165 106.100 114.135 ;
        RECT 119.285 111.735 119.710 117.130 ;
        RECT 120.330 116.620 121.330 116.790 ;
        RECT 120.100 112.410 120.270 116.450 ;
        RECT 121.390 112.410 121.560 116.450 ;
        RECT 121.950 114.735 122.670 117.130 ;
        RECT 123.290 116.620 124.290 116.790 ;
        RECT 123.060 115.410 123.230 116.450 ;
        RECT 124.350 115.410 124.520 116.450 ;
        RECT 123.290 115.070 124.290 115.240 ;
        RECT 124.900 114.735 125.370 117.130 ;
        RECT 120.330 112.070 121.330 112.240 ;
        RECT 121.950 111.735 125.370 114.735 ;
        RECT 119.285 111.210 125.370 111.735 ;
        RECT 101.160 110.425 104.175 111.165 ;
        RECT 104.790 110.660 105.290 110.830 ;
        RECT 104.560 110.425 104.730 110.445 ;
        RECT 101.160 109.925 104.760 110.425 ;
        RECT 101.160 109.180 104.175 109.925 ;
        RECT 104.560 109.905 104.730 109.925 ;
        RECT 105.350 109.905 105.520 110.445 ;
        RECT 104.790 109.520 105.290 109.690 ;
        RECT 105.920 109.180 106.090 111.165 ;
        RECT 98.540 109.005 100.540 109.175 ;
        RECT 101.160 109.010 106.090 109.180 ;
        RECT 101.160 109.000 104.175 109.010 ;
        RECT 101.160 108.665 102.070 109.000 ;
        RECT 97.740 108.495 102.070 108.665 ;
        RECT 81.750 108.480 82.585 108.490 ;
        RECT 101.160 108.480 102.070 108.495 ;
        RECT 79.625 107.470 80.295 107.480 ;
        RECT 79.625 107.300 86.000 107.470 ;
        RECT 103.440 107.465 104.185 107.475 ;
        RECT 79.625 106.545 80.295 107.300 ;
        RECT 80.910 106.790 82.910 106.960 ;
        RECT 83.200 106.790 85.200 106.960 ;
        RECT 80.680 106.545 80.850 106.620 ;
        RECT 79.625 102.655 80.855 106.545 ;
        RECT 79.625 101.915 80.295 102.655 ;
        RECT 80.680 102.580 80.850 102.655 ;
        RECT 82.970 102.580 83.140 106.620 ;
        RECT 85.260 105.485 85.430 106.620 ;
        RECT 85.830 105.485 86.000 107.300 ;
        RECT 97.740 107.295 106.090 107.465 ;
        RECT 97.740 105.485 97.910 107.295 ;
        RECT 98.540 106.785 100.540 106.955 ;
        RECT 100.830 106.785 102.830 106.955 ;
        RECT 98.310 105.485 98.480 106.615 ;
        RECT 85.255 105.470 86.540 105.485 ;
        RECT 97.190 105.470 98.485 105.485 ;
        RECT 85.255 105.300 98.485 105.470 ;
        RECT 85.255 102.655 86.540 105.300 ;
        RECT 87.150 104.790 91.150 104.960 ;
        RECT 85.260 102.580 85.430 102.655 ;
        RECT 80.910 102.240 82.910 102.410 ;
        RECT 83.200 102.240 85.200 102.410 ;
        RECT 85.810 101.915 86.540 102.655 ;
        RECT 86.920 102.580 87.090 104.620 ;
        RECT 91.210 102.580 91.380 104.620 ;
        RECT 87.150 102.240 91.150 102.410 ;
        RECT 91.780 101.915 91.950 105.300 ;
        RECT 92.580 104.790 96.580 104.960 ;
        RECT 92.350 102.580 92.520 104.620 ;
        RECT 96.640 102.580 96.810 104.620 ;
        RECT 97.190 102.650 98.485 105.300 ;
        RECT 92.580 102.240 96.580 102.410 ;
        RECT 97.190 101.915 97.920 102.650 ;
        RECT 98.310 102.575 98.480 102.650 ;
        RECT 100.600 102.575 100.770 106.615 ;
        RECT 102.890 106.540 103.060 106.615 ;
        RECT 103.440 106.595 104.185 107.295 ;
        RECT 104.790 106.785 105.290 106.955 ;
        RECT 104.560 106.595 104.730 106.615 ;
        RECT 103.440 106.540 104.760 106.595 ;
        RECT 102.885 104.795 104.760 106.540 ;
        RECT 102.885 104.110 104.185 104.795 ;
        RECT 104.560 104.775 104.730 104.795 ;
        RECT 105.350 104.775 105.520 106.615 ;
        RECT 104.790 104.435 105.290 104.605 ;
        RECT 105.920 104.110 106.090 107.295 ;
        RECT 102.885 102.650 106.120 104.110 ;
        RECT 102.890 102.575 103.060 102.650 ;
        RECT 98.540 102.235 100.540 102.405 ;
        RECT 100.830 102.235 102.830 102.405 ;
        RECT 103.445 101.915 106.120 102.650 ;
        RECT 79.625 100.505 106.120 101.915 ;
        RECT 79.625 99.995 106.125 100.505 ;
      LAYER met1 ;
        RECT 77.700 176.000 78.300 217.900 ;
        RECT 90.850 197.240 120.290 197.720 ;
        RECT 92.300 196.840 92.620 197.100 ;
        RECT 93.235 196.175 93.525 196.405 ;
        RECT 94.615 196.175 94.905 196.405 ;
        RECT 93.310 195.680 93.450 196.175 ;
        RECT 94.690 196.020 94.830 196.175 ;
        RECT 95.520 196.160 95.840 196.420 ;
        RECT 101.040 196.020 101.360 196.080 ;
        RECT 94.690 195.880 101.360 196.020 ;
        RECT 101.040 195.820 101.360 195.880 ;
        RECT 105.640 195.680 105.960 195.740 ;
        RECT 93.310 195.540 105.960 195.680 ;
        RECT 105.640 195.480 105.960 195.540 ;
        RECT 93.680 195.140 94.000 195.400 ;
        RECT 96.455 195.340 96.745 195.385 ;
        RECT 100.580 195.340 100.900 195.400 ;
        RECT 96.455 195.200 100.900 195.340 ;
        RECT 96.455 195.155 96.745 195.200 ;
        RECT 100.580 195.140 100.900 195.200 ;
        RECT 90.850 194.520 120.290 195.000 ;
        RECT 108.860 192.960 109.180 193.020 ;
        RECT 109.795 192.960 110.085 193.005 ;
        RECT 108.860 192.820 110.085 192.960 ;
        RECT 108.860 192.760 109.180 192.820 ;
        RECT 109.795 192.775 110.085 192.820 ;
        RECT 116.220 192.420 116.540 192.680 ;
        RECT 90.850 191.800 120.290 192.280 ;
        RECT 98.760 191.260 99.050 191.305 ;
        RECT 100.580 191.260 100.870 191.305 ;
        RECT 98.760 191.120 100.870 191.260 ;
        RECT 98.760 191.075 99.050 191.120 ;
        RECT 100.580 191.075 100.870 191.120 ;
        RECT 101.520 191.260 101.810 191.305 ;
        RECT 104.720 191.260 105.040 191.320 ;
        RECT 105.200 191.260 105.490 191.305 ;
        RECT 101.520 191.120 105.490 191.260 ;
        RECT 101.520 191.075 101.810 191.120 ;
        RECT 100.675 190.920 100.870 191.075 ;
        RECT 104.720 191.060 105.040 191.120 ;
        RECT 105.200 191.075 105.490 191.120 ;
        RECT 103.820 190.920 104.110 190.965 ;
        RECT 100.675 190.780 104.110 190.920 ;
        RECT 103.820 190.735 104.110 190.780 ;
        RECT 107.035 190.735 107.325 190.965 ;
        RECT 97.835 190.580 98.125 190.625 ;
        RECT 99.660 190.580 99.980 190.640 ;
        RECT 97.835 190.440 99.980 190.580 ;
        RECT 97.835 190.395 98.125 190.440 ;
        RECT 99.660 190.380 99.980 190.440 ;
        RECT 103.360 190.580 103.650 190.625 ;
        RECT 106.580 190.580 106.870 190.625 ;
        RECT 103.360 190.440 106.870 190.580 ;
        RECT 103.360 190.395 103.650 190.440 ;
        RECT 106.580 190.395 106.870 190.440 ;
        RECT 98.300 190.240 98.590 190.285 ;
        RECT 100.140 190.240 100.430 190.285 ;
        RECT 103.820 190.240 104.110 190.285 ;
        RECT 98.300 190.100 104.110 190.240 ;
        RECT 98.300 190.055 98.590 190.100 ;
        RECT 100.140 190.055 100.430 190.100 ;
        RECT 103.820 190.055 104.110 190.100 ;
        RECT 105.180 190.240 105.500 190.300 ;
        RECT 107.110 190.240 107.250 190.735 ;
        RECT 105.180 190.100 107.250 190.240 ;
        RECT 105.180 190.040 105.500 190.100 ;
        RECT 109.335 189.900 109.625 189.945 ;
        RECT 112.540 189.900 112.860 189.960 ;
        RECT 109.335 189.760 112.860 189.900 ;
        RECT 109.335 189.715 109.625 189.760 ;
        RECT 112.540 189.700 112.860 189.760 ;
        RECT 90.850 189.080 120.290 189.560 ;
        RECT 100.580 188.880 100.900 188.940 ;
        RECT 104.275 188.880 104.565 188.925 ;
        RECT 104.720 188.880 105.040 188.940 ;
        RECT 100.580 188.740 101.270 188.880 ;
        RECT 100.580 188.680 100.900 188.740 ;
        RECT 94.105 188.540 94.395 188.585 ;
        RECT 95.995 188.540 96.285 188.585 ;
        RECT 99.115 188.540 99.405 188.585 ;
        RECT 94.105 188.400 99.405 188.540 ;
        RECT 94.105 188.355 94.395 188.400 ;
        RECT 95.995 188.355 96.285 188.400 ;
        RECT 99.115 188.355 99.405 188.400 ;
        RECT 94.615 188.200 94.905 188.245 ;
        RECT 100.580 188.200 100.900 188.260 ;
        RECT 94.615 188.060 100.900 188.200 ;
        RECT 94.615 188.015 94.905 188.060 ;
        RECT 100.580 188.000 100.900 188.060 ;
        RECT 93.220 187.660 93.540 187.920 ;
        RECT 93.700 187.860 93.990 187.905 ;
        RECT 95.535 187.860 95.825 187.905 ;
        RECT 99.115 187.860 99.405 187.905 ;
        RECT 93.700 187.720 99.405 187.860 ;
        RECT 93.700 187.675 93.990 187.720 ;
        RECT 95.535 187.675 95.825 187.720 ;
        RECT 99.115 187.675 99.405 187.720 ;
        RECT 100.195 187.565 100.485 187.880 ;
        RECT 96.895 187.520 97.545 187.565 ;
        RECT 100.195 187.520 100.785 187.565 ;
        RECT 101.130 187.520 101.270 188.740 ;
        RECT 104.275 188.740 105.040 188.880 ;
        RECT 104.275 188.695 104.565 188.740 ;
        RECT 104.720 188.680 105.040 188.740 ;
        RECT 105.640 188.925 105.960 188.940 ;
        RECT 105.640 188.695 106.175 188.925 ;
        RECT 105.640 188.680 105.960 188.695 ;
        RECT 108.515 188.540 108.805 188.585 ;
        RECT 111.635 188.540 111.925 188.585 ;
        RECT 113.525 188.540 113.815 188.585 ;
        RECT 108.515 188.400 113.815 188.540 ;
        RECT 108.515 188.355 108.805 188.400 ;
        RECT 111.635 188.355 111.925 188.400 ;
        RECT 113.525 188.355 113.815 188.400 ;
        RECT 101.745 188.200 102.035 188.245 ;
        RECT 113.015 188.200 113.305 188.245 ;
        RECT 101.745 188.060 113.305 188.200 ;
        RECT 101.745 188.015 102.035 188.060 ;
        RECT 113.015 188.015 113.305 188.060 ;
        RECT 114.395 188.200 114.685 188.245 ;
        RECT 116.220 188.200 116.540 188.260 ;
        RECT 114.395 188.060 116.540 188.200 ;
        RECT 114.395 188.015 114.685 188.060 ;
        RECT 116.220 188.000 116.540 188.060 ;
        RECT 101.960 187.520 102.280 187.580 ;
        RECT 96.895 187.380 102.280 187.520 ;
        RECT 96.895 187.335 97.545 187.380 ;
        RECT 100.495 187.335 100.785 187.380 ;
        RECT 101.960 187.320 102.280 187.380 ;
        RECT 103.355 187.520 103.645 187.565 ;
        RECT 105.180 187.520 105.500 187.580 ;
        RECT 103.355 187.380 105.500 187.520 ;
        RECT 103.355 187.335 103.645 187.380 ;
        RECT 105.180 187.320 105.500 187.380 ;
        RECT 105.640 187.520 105.960 187.580 ;
        RECT 107.435 187.565 107.725 187.880 ;
        RECT 108.515 187.860 108.805 187.905 ;
        RECT 112.095 187.860 112.385 187.905 ;
        RECT 113.930 187.860 114.220 187.905 ;
        RECT 108.515 187.720 114.220 187.860 ;
        RECT 108.515 187.675 108.805 187.720 ;
        RECT 112.095 187.675 112.385 187.720 ;
        RECT 113.930 187.675 114.220 187.720 ;
        RECT 107.135 187.520 107.725 187.565 ;
        RECT 110.375 187.520 111.025 187.565 ;
        RECT 105.640 187.380 111.025 187.520 ;
        RECT 105.640 187.320 105.960 187.380 ;
        RECT 107.135 187.335 107.425 187.380 ;
        RECT 110.375 187.335 111.025 187.380 ;
        RECT 99.660 187.180 99.980 187.240 ;
        RECT 104.720 187.180 105.040 187.240 ;
        RECT 99.660 187.040 105.040 187.180 ;
        RECT 99.660 186.980 99.980 187.040 ;
        RECT 104.720 186.980 105.040 187.040 ;
        RECT 90.850 186.360 120.290 186.840 ;
        RECT 101.040 185.960 101.360 186.220 ;
        RECT 105.210 185.865 105.470 185.910 ;
        RECT 105.190 185.820 105.480 185.865 ;
        RECT 108.870 185.820 109.160 185.865 ;
        RECT 105.190 185.680 109.160 185.820 ;
        RECT 105.190 185.635 105.480 185.680 ;
        RECT 108.870 185.635 109.160 185.680 ;
        RECT 109.810 185.820 110.100 185.865 ;
        RECT 111.630 185.820 111.920 185.865 ;
        RECT 109.810 185.680 111.920 185.820 ;
        RECT 109.810 185.635 110.100 185.680 ;
        RECT 111.630 185.635 111.920 185.680 ;
        RECT 105.210 185.590 105.470 185.635 ;
        RECT 93.235 185.480 93.525 185.525 ;
        RECT 97.360 185.480 97.680 185.540 ;
        RECT 93.235 185.340 97.680 185.480 ;
        RECT 93.235 185.295 93.525 185.340 ;
        RECT 97.360 185.280 97.680 185.340 ;
        RECT 101.960 185.480 102.280 185.540 ;
        RECT 103.355 185.480 103.645 185.525 ;
        RECT 101.960 185.340 103.645 185.480 ;
        RECT 101.960 185.280 102.280 185.340 ;
        RECT 103.355 185.295 103.645 185.340 ;
        RECT 106.570 185.480 106.860 185.525 ;
        RECT 109.810 185.480 110.005 185.635 ;
        RECT 106.570 185.340 110.005 185.480 ;
        RECT 106.570 185.295 106.860 185.340 ;
        RECT 103.430 184.800 103.570 185.295 ;
        RECT 112.540 185.280 112.860 185.540 ;
        RECT 118.535 185.480 118.825 185.525 ;
        RECT 119.900 185.480 120.220 185.540 ;
        RECT 118.535 185.340 120.220 185.480 ;
        RECT 118.535 185.295 118.825 185.340 ;
        RECT 119.900 185.280 120.220 185.340 ;
        RECT 103.810 185.140 104.100 185.185 ;
        RECT 107.030 185.140 107.320 185.185 ;
        RECT 103.810 185.000 107.320 185.140 ;
        RECT 103.810 184.955 104.100 185.000 ;
        RECT 107.030 184.955 107.320 185.000 ;
        RECT 108.400 185.140 108.720 185.200 ;
        RECT 110.715 185.140 111.005 185.185 ;
        RECT 108.400 185.000 112.770 185.140 ;
        RECT 108.400 184.940 108.720 185.000 ;
        RECT 110.715 184.955 111.005 185.000 ;
        RECT 112.630 184.860 112.770 185.000 ;
        RECT 105.640 184.800 105.960 184.860 ;
        RECT 103.430 184.660 105.960 184.800 ;
        RECT 105.640 184.600 105.960 184.660 ;
        RECT 106.570 184.800 106.860 184.845 ;
        RECT 110.250 184.800 110.540 184.845 ;
        RECT 112.090 184.800 112.380 184.845 ;
        RECT 106.570 184.660 112.380 184.800 ;
        RECT 106.570 184.615 106.860 184.660 ;
        RECT 110.250 184.615 110.540 184.660 ;
        RECT 112.090 184.615 112.380 184.660 ;
        RECT 112.540 184.800 112.860 184.860 ;
        RECT 117.615 184.800 117.905 184.845 ;
        RECT 112.540 184.660 117.905 184.800 ;
        RECT 112.540 184.600 112.860 184.660 ;
        RECT 117.615 184.615 117.905 184.660 ;
        RECT 89.540 184.460 89.860 184.520 ;
        RECT 92.315 184.460 92.605 184.505 ;
        RECT 89.540 184.320 92.605 184.460 ;
        RECT 89.540 184.260 89.860 184.320 ;
        RECT 92.315 184.275 92.605 184.320 ;
        RECT 90.850 183.640 120.290 184.120 ;
        RECT 97.360 183.440 97.680 183.500 ;
        RECT 97.360 183.300 115.990 183.440 ;
        RECT 97.360 183.240 97.680 183.300 ;
        RECT 94.105 183.100 94.395 183.145 ;
        RECT 95.995 183.100 96.285 183.145 ;
        RECT 99.115 183.100 99.405 183.145 ;
        RECT 94.105 182.960 99.405 183.100 ;
        RECT 94.105 182.915 94.395 182.960 ;
        RECT 95.995 182.915 96.285 182.960 ;
        RECT 99.115 182.915 99.405 182.960 ;
        RECT 109.790 183.100 110.080 183.145 ;
        RECT 113.470 183.100 113.760 183.145 ;
        RECT 115.310 183.100 115.600 183.145 ;
        RECT 109.790 182.960 115.600 183.100 ;
        RECT 109.790 182.915 110.080 182.960 ;
        RECT 113.470 182.915 113.760 182.960 ;
        RECT 115.310 182.915 115.600 182.960 ;
        RECT 94.615 182.760 94.905 182.805 ;
        RECT 104.720 182.760 105.040 182.820 ;
        RECT 94.615 182.620 105.040 182.760 ;
        RECT 94.615 182.575 94.905 182.620 ;
        RECT 104.720 182.560 105.040 182.620 ;
        RECT 107.030 182.760 107.320 182.805 ;
        RECT 110.250 182.760 110.540 182.805 ;
        RECT 107.030 182.620 110.540 182.760 ;
        RECT 107.030 182.575 107.320 182.620 ;
        RECT 110.250 182.575 110.540 182.620 ;
        RECT 112.540 182.760 112.860 182.820 ;
        RECT 115.850 182.805 115.990 183.300 ;
        RECT 113.935 182.760 114.225 182.805 ;
        RECT 112.540 182.620 114.225 182.760 ;
        RECT 112.540 182.560 112.860 182.620 ;
        RECT 113.935 182.575 114.225 182.620 ;
        RECT 115.775 182.575 116.065 182.805 ;
        RECT 93.220 182.220 93.540 182.480 ;
        RECT 93.700 182.420 93.990 182.465 ;
        RECT 95.535 182.420 95.825 182.465 ;
        RECT 99.115 182.420 99.405 182.465 ;
        RECT 93.700 182.280 99.405 182.420 ;
        RECT 93.700 182.235 93.990 182.280 ;
        RECT 95.535 182.235 95.825 182.280 ;
        RECT 99.115 182.235 99.405 182.280 ;
        RECT 96.895 182.080 97.545 182.125 ;
        RECT 97.820 182.080 98.140 182.140 ;
        RECT 100.195 182.125 100.485 182.440 ;
        RECT 101.040 182.420 101.360 182.480 ;
        RECT 101.745 182.420 102.035 182.465 ;
        RECT 101.040 182.280 102.035 182.420 ;
        RECT 101.040 182.220 101.360 182.280 ;
        RECT 101.745 182.235 102.035 182.280 ;
        RECT 104.260 182.420 104.580 182.480 ;
        RECT 105.640 182.420 105.960 182.480 ;
        RECT 106.575 182.420 106.865 182.465 ;
        RECT 104.260 182.280 106.865 182.420 ;
        RECT 104.260 182.220 104.580 182.280 ;
        RECT 105.640 182.220 105.960 182.280 ;
        RECT 106.575 182.235 106.865 182.280 ;
        RECT 109.790 182.420 110.080 182.465 ;
        RECT 109.790 182.280 113.225 182.420 ;
        RECT 109.790 182.235 110.080 182.280 ;
        RECT 113.030 182.125 113.225 182.280 ;
        RECT 100.195 182.080 100.785 182.125 ;
        RECT 96.895 181.940 100.785 182.080 ;
        RECT 96.895 181.895 97.545 181.940 ;
        RECT 97.820 181.880 98.140 181.940 ;
        RECT 100.495 181.895 100.785 181.940 ;
        RECT 103.355 182.080 103.645 182.125 ;
        RECT 108.410 182.080 108.700 182.125 ;
        RECT 112.090 182.080 112.380 182.125 ;
        RECT 103.355 181.940 112.380 182.080 ;
        RECT 103.355 181.895 103.645 181.940 ;
        RECT 108.410 181.895 108.700 181.940 ;
        RECT 112.090 181.895 112.380 181.940 ;
        RECT 113.030 182.080 113.320 182.125 ;
        RECT 114.850 182.080 115.140 182.125 ;
        RECT 113.030 181.940 115.140 182.080 ;
        RECT 113.030 181.895 113.320 181.940 ;
        RECT 114.850 181.895 115.140 181.940 ;
        RECT 104.275 181.740 104.565 181.785 ;
        RECT 105.640 181.740 105.960 181.800 ;
        RECT 104.275 181.600 105.960 181.740 ;
        RECT 104.275 181.555 104.565 181.600 ;
        RECT 105.640 181.540 105.960 181.600 ;
        RECT 90.850 180.920 120.290 181.400 ;
        RECT 96.915 180.720 97.205 180.765 ;
        RECT 97.360 180.720 97.680 180.780 ;
        RECT 96.915 180.580 97.680 180.720 ;
        RECT 96.915 180.535 97.205 180.580 ;
        RECT 97.360 180.520 97.680 180.580 ;
        RECT 101.500 180.720 101.820 180.780 ;
        RECT 101.500 180.580 108.630 180.720 ;
        RECT 101.500 180.520 101.820 180.580 ;
        RECT 101.050 180.380 101.340 180.425 ;
        RECT 101.960 180.380 102.280 180.440 ;
        RECT 104.730 180.380 105.020 180.425 ;
        RECT 101.050 180.240 105.020 180.380 ;
        RECT 101.050 180.195 101.340 180.240 ;
        RECT 101.960 180.180 102.280 180.240 ;
        RECT 104.730 180.195 105.020 180.240 ;
        RECT 105.670 180.380 105.960 180.425 ;
        RECT 107.490 180.380 107.780 180.425 ;
        RECT 105.670 180.240 107.780 180.380 ;
        RECT 105.670 180.195 105.960 180.240 ;
        RECT 107.490 180.195 107.780 180.240 ;
        RECT 97.820 180.040 98.140 180.100 ;
        RECT 99.215 180.040 99.505 180.085 ;
        RECT 101.500 180.040 101.820 180.100 ;
        RECT 97.820 179.900 101.820 180.040 ;
        RECT 97.820 179.840 98.140 179.900 ;
        RECT 99.215 179.855 99.505 179.900 ;
        RECT 101.500 179.840 101.820 179.900 ;
        RECT 102.430 180.040 102.720 180.085 ;
        RECT 105.670 180.040 105.865 180.195 ;
        RECT 102.430 179.900 105.865 180.040 ;
        RECT 106.575 180.040 106.865 180.085 ;
        RECT 107.940 180.040 108.260 180.100 ;
        RECT 108.490 180.085 108.630 180.580 ;
        RECT 106.575 179.900 108.260 180.040 ;
        RECT 102.430 179.855 102.720 179.900 ;
        RECT 106.575 179.855 106.865 179.900 ;
        RECT 107.940 179.840 108.260 179.900 ;
        RECT 108.415 179.855 108.705 180.085 ;
        RECT 99.670 179.700 99.960 179.745 ;
        RECT 102.890 179.700 103.180 179.745 ;
        RECT 99.670 179.560 103.180 179.700 ;
        RECT 99.670 179.515 99.960 179.560 ;
        RECT 102.890 179.515 103.180 179.560 ;
        RECT 102.430 179.360 102.720 179.405 ;
        RECT 106.110 179.360 106.400 179.405 ;
        RECT 107.950 179.360 108.240 179.405 ;
        RECT 102.430 179.220 108.240 179.360 ;
        RECT 102.430 179.175 102.720 179.220 ;
        RECT 106.110 179.175 106.400 179.220 ;
        RECT 107.950 179.175 108.240 179.220 ;
        RECT 101.500 179.020 101.820 179.080 ;
        RECT 104.260 179.020 104.580 179.080 ;
        RECT 101.500 178.880 104.580 179.020 ;
        RECT 101.500 178.820 101.820 178.880 ;
        RECT 104.260 178.820 104.580 178.880 ;
        RECT 90.850 178.200 120.290 178.680 ;
        RECT 104.720 177.800 105.040 178.060 ;
        RECT 94.105 177.660 94.395 177.705 ;
        RECT 95.995 177.660 96.285 177.705 ;
        RECT 99.115 177.660 99.405 177.705 ;
        RECT 94.105 177.520 99.405 177.660 ;
        RECT 94.105 177.475 94.395 177.520 ;
        RECT 95.995 177.475 96.285 177.520 ;
        RECT 99.115 177.475 99.405 177.520 ;
        RECT 100.580 177.660 100.900 177.720 ;
        RECT 101.745 177.660 102.035 177.705 ;
        RECT 100.580 177.520 102.035 177.660 ;
        RECT 100.580 177.460 100.900 177.520 ;
        RECT 101.745 177.475 102.035 177.520 ;
        RECT 109.335 177.660 109.625 177.705 ;
        RECT 112.095 177.660 112.385 177.705 ;
        RECT 113.895 177.660 114.185 177.705 ;
        RECT 109.335 177.520 114.185 177.660 ;
        RECT 109.335 177.475 109.625 177.520 ;
        RECT 112.095 177.475 112.385 177.520 ;
        RECT 113.895 177.475 114.185 177.520 ;
        RECT 94.615 177.320 94.905 177.365 ;
        RECT 101.040 177.320 101.360 177.380 ;
        RECT 94.615 177.180 101.360 177.320 ;
        RECT 94.615 177.135 94.905 177.180 ;
        RECT 101.040 177.120 101.360 177.180 ;
        RECT 104.720 177.320 105.040 177.380 ;
        RECT 112.555 177.320 112.845 177.365 ;
        RECT 104.720 177.180 112.845 177.320 ;
        RECT 104.720 177.120 105.040 177.180 ;
        RECT 112.555 177.135 112.845 177.180 ;
        RECT 114.395 177.320 114.685 177.365 ;
        RECT 116.220 177.320 116.540 177.380 ;
        RECT 114.395 177.180 116.540 177.320 ;
        RECT 114.395 177.135 114.685 177.180 ;
        RECT 116.220 177.120 116.540 177.180 ;
        RECT 93.220 176.780 93.540 177.040 ;
        RECT 93.700 176.980 93.990 177.025 ;
        RECT 95.535 176.980 95.825 177.025 ;
        RECT 99.115 176.980 99.405 177.025 ;
        RECT 93.700 176.840 99.405 176.980 ;
        RECT 93.700 176.795 93.990 176.840 ;
        RECT 95.535 176.795 95.825 176.840 ;
        RECT 99.115 176.795 99.405 176.840 ;
        RECT 100.195 176.685 100.485 177.000 ;
        RECT 101.960 176.980 102.280 177.040 ;
        RECT 103.355 176.980 103.645 177.025 ;
        RECT 101.960 176.840 103.645 176.980 ;
        RECT 101.960 176.780 102.280 176.840 ;
        RECT 103.355 176.795 103.645 176.840 ;
        RECT 109.295 176.980 109.585 177.025 ;
        RECT 109.295 176.840 111.850 176.980 ;
        RECT 109.295 176.795 109.585 176.840 ;
        RECT 96.895 176.640 97.545 176.685 ;
        RECT 100.195 176.640 100.785 176.685 ;
        RECT 101.500 176.640 101.820 176.700 ;
        RECT 111.635 176.685 111.850 176.840 ;
        RECT 107.495 176.640 107.785 176.685 ;
        RECT 110.715 176.640 111.005 176.685 ;
        RECT 96.895 176.500 111.005 176.640 ;
        RECT 96.895 176.455 97.545 176.500 ;
        RECT 100.495 176.455 100.785 176.500 ;
        RECT 101.500 176.440 101.820 176.500 ;
        RECT 107.495 176.455 107.785 176.500 ;
        RECT 110.715 176.455 111.005 176.500 ;
        RECT 111.635 176.640 111.925 176.685 ;
        RECT 113.475 176.640 113.765 176.685 ;
        RECT 111.635 176.500 113.765 176.640 ;
        RECT 111.635 176.455 111.925 176.500 ;
        RECT 113.475 176.455 113.765 176.500 ;
        RECT 105.180 176.300 105.500 176.360 ;
        RECT 106.115 176.300 106.405 176.345 ;
        RECT 105.180 176.160 106.405 176.300 ;
        RECT 105.180 176.100 105.500 176.160 ;
        RECT 106.115 176.115 106.405 176.160 ;
        RECT 90.850 175.480 120.290 175.960 ;
        RECT 105.180 175.280 105.500 175.340 ;
        RECT 104.350 175.140 105.500 175.280 ;
        RECT 100.130 174.940 100.420 174.985 ;
        RECT 103.810 174.940 104.100 174.985 ;
        RECT 104.350 174.940 104.490 175.140 ;
        RECT 105.180 175.080 105.500 175.140 ;
        RECT 100.130 174.800 104.490 174.940 ;
        RECT 104.750 174.940 105.040 174.985 ;
        RECT 106.570 174.940 106.860 174.985 ;
        RECT 104.750 174.800 106.860 174.940 ;
        RECT 100.130 174.755 100.420 174.800 ;
        RECT 103.810 174.755 104.100 174.800 ;
        RECT 104.750 174.755 105.040 174.800 ;
        RECT 106.570 174.755 106.860 174.800 ;
        RECT 93.235 174.415 93.525 174.645 ;
        RECT 94.615 174.415 94.905 174.645 ;
        RECT 98.295 174.600 98.585 174.645 ;
        RECT 101.040 174.600 101.360 174.660 ;
        RECT 98.295 174.460 101.360 174.600 ;
        RECT 98.295 174.415 98.585 174.460 ;
        RECT 89.540 173.920 89.860 173.980 ;
        RECT 92.315 173.920 92.605 173.965 ;
        RECT 89.540 173.780 92.605 173.920 ;
        RECT 93.310 173.920 93.450 174.415 ;
        RECT 94.690 174.260 94.830 174.415 ;
        RECT 101.040 174.400 101.360 174.460 ;
        RECT 101.510 174.600 101.800 174.645 ;
        RECT 104.750 174.600 104.945 174.755 ;
        RECT 101.510 174.460 104.945 174.600 ;
        RECT 105.655 174.600 105.945 174.645 ;
        RECT 108.400 174.600 108.720 174.660 ;
        RECT 105.655 174.460 108.720 174.600 ;
        RECT 101.510 174.415 101.800 174.460 ;
        RECT 105.655 174.415 105.945 174.460 ;
        RECT 108.400 174.400 108.720 174.460 ;
        RECT 95.995 174.260 96.285 174.305 ;
        RECT 94.690 174.120 96.285 174.260 ;
        RECT 95.995 174.075 96.285 174.120 ;
        RECT 98.750 174.260 99.040 174.305 ;
        RECT 101.970 174.260 102.260 174.305 ;
        RECT 98.750 174.120 102.260 174.260 ;
        RECT 98.750 174.075 99.040 174.120 ;
        RECT 101.970 174.075 102.260 174.120 ;
        RECT 107.495 174.075 107.785 174.305 ;
        RECT 101.510 173.920 101.800 173.965 ;
        RECT 105.190 173.920 105.480 173.965 ;
        RECT 107.030 173.920 107.320 173.965 ;
        RECT 93.310 173.780 101.270 173.920 ;
        RECT 89.540 173.720 89.860 173.780 ;
        RECT 92.315 173.735 92.605 173.780 ;
        RECT 93.680 173.380 94.000 173.640 ;
        RECT 101.130 173.580 101.270 173.780 ;
        RECT 101.510 173.780 107.320 173.920 ;
        RECT 101.510 173.735 101.800 173.780 ;
        RECT 105.190 173.735 105.480 173.780 ;
        RECT 107.030 173.735 107.320 173.780 ;
        RECT 105.640 173.580 105.960 173.640 ;
        RECT 107.570 173.580 107.710 174.075 ;
        RECT 101.130 173.440 107.710 173.580 ;
        RECT 105.640 173.380 105.960 173.440 ;
        RECT 90.850 172.760 120.290 173.240 ;
        RECT 93.220 172.560 93.540 172.620 ;
        RECT 93.695 172.560 93.985 172.605 ;
        RECT 93.220 172.420 93.985 172.560 ;
        RECT 93.220 172.360 93.540 172.420 ;
        RECT 93.695 172.375 93.985 172.420 ;
        RECT 102.435 172.560 102.725 172.605 ;
        RECT 104.720 172.560 105.040 172.620 ;
        RECT 102.435 172.420 105.040 172.560 ;
        RECT 102.435 172.375 102.725 172.420 ;
        RECT 104.720 172.360 105.040 172.420 ;
        RECT 106.575 172.560 106.865 172.605 ;
        RECT 108.860 172.560 109.180 172.620 ;
        RECT 106.575 172.420 109.180 172.560 ;
        RECT 106.575 172.375 106.865 172.420 ;
        RECT 106.650 171.880 106.790 172.375 ;
        RECT 108.860 172.360 109.180 172.420 ;
        RECT 101.130 171.740 106.790 171.880 ;
        RECT 101.130 171.585 101.270 171.740 ;
        RECT 101.055 171.355 101.345 171.585 ;
        RECT 103.355 171.540 103.645 171.585 ;
        RECT 105.180 171.540 105.500 171.600 ;
        RECT 103.355 171.400 105.500 171.540 ;
        RECT 103.355 171.355 103.645 171.400 ;
        RECT 105.180 171.340 105.500 171.400 ;
        RECT 113.000 171.340 113.320 171.600 ;
        RECT 90.850 170.040 120.290 170.520 ;
        RECT 47.600 153.320 48.500 157.100 ;
        RECT 47.565 146.800 48.565 153.320 ;
        RECT 58.195 152.800 59.195 153.335 ;
        RECT 61.100 153.295 62.100 157.100 ;
        RECT 49.790 152.475 51.645 152.595 ;
        RECT 55.075 152.475 56.925 152.600 ;
        RECT 49.715 152.245 51.715 152.475 ;
        RECT 55.000 152.245 57.000 152.475 ;
        RECT 58.145 152.435 59.195 152.800 ;
        RECT 49.790 152.235 51.645 152.245 ;
        RECT 55.075 152.240 56.925 152.245 ;
        RECT 49.325 151.865 49.555 152.195 ;
        RECT 51.875 151.865 52.105 152.195 ;
        RECT 52.850 151.865 53.810 151.895 ;
        RECT 54.565 151.865 54.795 152.195 ;
        RECT 57.205 151.865 57.435 152.195 ;
        RECT 49.325 151.565 57.435 151.865 ;
        RECT 49.325 151.235 49.555 151.565 ;
        RECT 51.875 151.235 52.105 151.565 ;
        RECT 52.850 151.535 53.810 151.565 ;
        RECT 54.565 151.235 54.795 151.565 ;
        RECT 57.205 151.235 57.435 151.565 ;
        RECT 49.715 150.955 51.715 151.185 ;
        RECT 55.000 150.955 57.000 151.185 ;
        RECT 49.770 150.815 51.660 150.955 ;
        RECT 55.055 150.815 56.945 150.955 ;
        RECT 49.770 150.615 56.945 150.815 ;
        RECT 49.790 150.045 51.640 150.175 ;
        RECT 49.715 149.815 51.715 150.045 ;
        RECT 49.325 149.675 49.555 149.765 ;
        RECT 51.875 149.675 52.105 149.765 ;
        RECT 53.420 149.675 53.820 150.615 ;
        RECT 55.075 150.045 56.920 150.180 ;
        RECT 55.000 149.815 57.000 150.045 ;
        RECT 54.565 149.675 54.795 149.765 ;
        RECT 57.205 149.675 57.435 149.765 ;
        RECT 49.325 149.465 57.435 149.675 ;
        RECT 49.325 149.395 49.645 149.465 ;
        RECT 51.785 149.395 54.935 149.465 ;
        RECT 57.070 149.395 57.435 149.465 ;
        RECT 49.325 149.305 49.555 149.395 ;
        RECT 49.790 149.255 51.640 149.320 ;
        RECT 51.875 149.305 52.105 149.395 ;
        RECT 49.715 149.025 51.715 149.255 ;
        RECT 49.325 148.885 49.555 148.975 ;
        RECT 49.790 148.960 51.640 149.025 ;
        RECT 51.875 148.885 52.105 148.975 ;
        RECT 53.420 148.885 53.820 149.395 ;
        RECT 54.565 149.305 54.795 149.395 ;
        RECT 55.080 149.255 56.925 149.320 ;
        RECT 57.205 149.305 57.435 149.395 ;
        RECT 55.000 149.025 57.000 149.255 ;
        RECT 54.565 148.885 54.795 148.975 ;
        RECT 55.080 148.960 56.925 149.025 ;
        RECT 57.205 148.885 57.435 148.975 ;
        RECT 49.325 148.815 49.645 148.885 ;
        RECT 51.785 148.815 54.935 148.885 ;
        RECT 57.070 148.815 57.435 148.885 ;
        RECT 49.325 148.675 57.435 148.815 ;
        RECT 49.325 148.605 49.645 148.675 ;
        RECT 51.785 148.605 54.935 148.675 ;
        RECT 57.070 148.605 57.435 148.675 ;
        RECT 49.325 148.515 49.555 148.605 ;
        RECT 49.795 148.465 51.640 148.530 ;
        RECT 51.875 148.515 52.105 148.605 ;
        RECT 49.715 148.235 51.715 148.465 ;
        RECT 49.325 148.095 49.555 148.185 ;
        RECT 49.795 148.170 51.640 148.235 ;
        RECT 51.875 148.095 52.105 148.185 ;
        RECT 53.420 148.095 53.820 148.605 ;
        RECT 54.565 148.515 54.795 148.605 ;
        RECT 55.090 148.465 56.940 148.530 ;
        RECT 57.205 148.515 57.435 148.605 ;
        RECT 55.000 148.235 57.000 148.465 ;
        RECT 54.565 148.095 54.795 148.185 ;
        RECT 55.090 148.170 56.940 148.235 ;
        RECT 57.205 148.095 57.435 148.185 ;
        RECT 49.325 148.025 49.645 148.095 ;
        RECT 51.785 148.025 54.935 148.095 ;
        RECT 57.070 148.025 57.435 148.095 ;
        RECT 49.325 147.885 57.435 148.025 ;
        RECT 49.325 147.815 49.650 147.885 ;
        RECT 51.785 147.815 54.935 147.885 ;
        RECT 57.070 147.815 57.435 147.885 ;
        RECT 49.325 147.725 49.555 147.815 ;
        RECT 49.795 147.675 51.640 147.740 ;
        RECT 51.875 147.725 52.105 147.815 ;
        RECT 49.715 147.445 51.715 147.675 ;
        RECT 49.795 147.380 51.640 147.445 ;
        RECT 54.100 147.305 54.360 147.815 ;
        RECT 54.565 147.725 54.795 147.815 ;
        RECT 55.090 147.675 56.915 147.740 ;
        RECT 57.205 147.725 57.435 147.815 ;
        RECT 55.000 147.445 57.000 147.675 ;
        RECT 54.565 147.305 54.795 147.395 ;
        RECT 55.090 147.380 56.915 147.445 ;
        RECT 57.205 147.305 57.435 147.395 ;
        RECT 54.100 147.235 54.935 147.305 ;
        RECT 57.070 147.235 57.435 147.305 ;
        RECT 54.100 147.095 57.435 147.235 ;
        RECT 54.100 147.025 54.935 147.095 ;
        RECT 57.070 147.025 57.435 147.095 ;
        RECT 54.100 146.515 54.360 147.025 ;
        RECT 54.565 146.935 54.795 147.025 ;
        RECT 55.075 146.885 56.925 146.950 ;
        RECT 57.205 146.935 57.435 147.025 ;
        RECT 55.000 146.655 57.000 146.885 ;
        RECT 54.565 146.515 54.795 146.605 ;
        RECT 55.075 146.590 56.925 146.655 ;
        RECT 57.205 146.515 57.435 146.605 ;
        RECT 54.100 146.445 54.935 146.515 ;
        RECT 57.070 146.445 57.435 146.515 ;
        RECT 54.100 146.305 57.435 146.445 ;
        RECT 54.100 146.235 54.935 146.305 ;
        RECT 57.070 146.235 57.435 146.305 ;
        RECT 54.565 146.145 54.795 146.235 ;
        RECT 55.080 146.095 56.915 146.160 ;
        RECT 57.205 146.145 57.435 146.235 ;
        RECT 55.000 145.865 57.000 146.095 ;
        RECT 55.080 145.800 56.915 145.865 ;
        RECT 58.195 145.100 59.195 152.435 ;
        RECT 61.095 153.200 62.100 153.295 ;
        RECT 61.095 146.775 62.095 153.200 ;
        RECT 71.725 152.775 72.725 153.310 ;
        RECT 63.320 152.450 65.175 152.570 ;
        RECT 68.605 152.450 70.455 152.575 ;
        RECT 63.245 152.220 65.245 152.450 ;
        RECT 68.530 152.220 70.530 152.450 ;
        RECT 71.675 152.410 72.725 152.775 ;
        RECT 63.320 152.210 65.175 152.220 ;
        RECT 68.605 152.215 70.455 152.220 ;
        RECT 62.855 151.840 63.085 152.170 ;
        RECT 65.405 151.840 65.635 152.170 ;
        RECT 66.380 151.840 67.340 151.870 ;
        RECT 68.095 151.840 68.325 152.170 ;
        RECT 70.735 151.840 70.965 152.170 ;
        RECT 62.855 151.540 70.965 151.840 ;
        RECT 62.855 151.210 63.085 151.540 ;
        RECT 65.405 151.210 65.635 151.540 ;
        RECT 66.380 151.510 67.340 151.540 ;
        RECT 68.095 151.210 68.325 151.540 ;
        RECT 70.735 151.210 70.965 151.540 ;
        RECT 63.245 150.930 65.245 151.160 ;
        RECT 68.530 150.930 70.530 151.160 ;
        RECT 63.300 150.790 65.190 150.930 ;
        RECT 68.585 150.790 70.475 150.930 ;
        RECT 63.300 150.590 70.475 150.790 ;
        RECT 63.320 150.020 65.170 150.150 ;
        RECT 63.245 149.790 65.245 150.020 ;
        RECT 62.855 149.650 63.085 149.740 ;
        RECT 65.405 149.650 65.635 149.740 ;
        RECT 66.950 149.650 67.350 150.590 ;
        RECT 68.605 150.020 70.450 150.155 ;
        RECT 68.530 149.790 70.530 150.020 ;
        RECT 68.095 149.650 68.325 149.740 ;
        RECT 70.735 149.650 70.965 149.740 ;
        RECT 62.855 149.440 70.965 149.650 ;
        RECT 62.855 149.370 63.175 149.440 ;
        RECT 65.315 149.370 68.465 149.440 ;
        RECT 70.600 149.370 70.965 149.440 ;
        RECT 62.855 149.280 63.085 149.370 ;
        RECT 63.320 149.230 65.170 149.295 ;
        RECT 65.405 149.280 65.635 149.370 ;
        RECT 63.245 149.000 65.245 149.230 ;
        RECT 62.855 148.860 63.085 148.950 ;
        RECT 63.320 148.935 65.170 149.000 ;
        RECT 65.405 148.860 65.635 148.950 ;
        RECT 66.950 148.860 67.350 149.370 ;
        RECT 68.095 149.280 68.325 149.370 ;
        RECT 68.610 149.230 70.455 149.295 ;
        RECT 70.735 149.280 70.965 149.370 ;
        RECT 68.530 149.000 70.530 149.230 ;
        RECT 68.095 148.860 68.325 148.950 ;
        RECT 68.610 148.935 70.455 149.000 ;
        RECT 70.735 148.860 70.965 148.950 ;
        RECT 62.855 148.790 63.175 148.860 ;
        RECT 65.315 148.790 68.465 148.860 ;
        RECT 70.600 148.790 70.965 148.860 ;
        RECT 62.855 148.650 70.965 148.790 ;
        RECT 62.855 148.580 63.175 148.650 ;
        RECT 65.315 148.580 68.465 148.650 ;
        RECT 70.600 148.580 70.965 148.650 ;
        RECT 62.855 148.490 63.085 148.580 ;
        RECT 63.325 148.440 65.170 148.505 ;
        RECT 65.405 148.490 65.635 148.580 ;
        RECT 63.245 148.210 65.245 148.440 ;
        RECT 62.855 148.070 63.085 148.160 ;
        RECT 63.325 148.145 65.170 148.210 ;
        RECT 65.405 148.070 65.635 148.160 ;
        RECT 66.950 148.070 67.350 148.580 ;
        RECT 68.095 148.490 68.325 148.580 ;
        RECT 68.620 148.440 70.470 148.505 ;
        RECT 70.735 148.490 70.965 148.580 ;
        RECT 68.530 148.210 70.530 148.440 ;
        RECT 68.095 148.070 68.325 148.160 ;
        RECT 68.620 148.145 70.470 148.210 ;
        RECT 70.735 148.070 70.965 148.160 ;
        RECT 62.855 148.000 63.175 148.070 ;
        RECT 65.315 148.000 68.465 148.070 ;
        RECT 70.600 148.000 70.965 148.070 ;
        RECT 62.855 147.860 70.965 148.000 ;
        RECT 62.855 147.790 63.180 147.860 ;
        RECT 65.315 147.790 68.465 147.860 ;
        RECT 70.600 147.790 70.965 147.860 ;
        RECT 62.855 147.700 63.085 147.790 ;
        RECT 63.325 147.650 65.170 147.715 ;
        RECT 65.405 147.700 65.635 147.790 ;
        RECT 63.245 147.420 65.245 147.650 ;
        RECT 63.325 147.355 65.170 147.420 ;
        RECT 67.630 147.280 67.890 147.790 ;
        RECT 68.095 147.700 68.325 147.790 ;
        RECT 68.620 147.650 70.445 147.715 ;
        RECT 70.735 147.700 70.965 147.790 ;
        RECT 68.530 147.420 70.530 147.650 ;
        RECT 68.095 147.280 68.325 147.370 ;
        RECT 68.620 147.355 70.445 147.420 ;
        RECT 70.735 147.280 70.965 147.370 ;
        RECT 67.630 147.210 68.465 147.280 ;
        RECT 70.600 147.210 70.965 147.280 ;
        RECT 67.630 147.070 70.965 147.210 ;
        RECT 67.630 147.000 68.465 147.070 ;
        RECT 70.600 147.000 70.965 147.070 ;
        RECT 67.630 146.490 67.890 147.000 ;
        RECT 68.095 146.910 68.325 147.000 ;
        RECT 68.605 146.860 70.455 146.925 ;
        RECT 70.735 146.910 70.965 147.000 ;
        RECT 68.530 146.630 70.530 146.860 ;
        RECT 68.095 146.490 68.325 146.580 ;
        RECT 68.605 146.565 70.455 146.630 ;
        RECT 70.735 146.490 70.965 146.580 ;
        RECT 67.630 146.420 68.465 146.490 ;
        RECT 70.600 146.420 70.965 146.490 ;
        RECT 67.630 146.280 70.965 146.420 ;
        RECT 67.630 146.210 68.465 146.280 ;
        RECT 70.600 146.210 70.965 146.280 ;
        RECT 68.095 146.120 68.325 146.210 ;
        RECT 68.610 146.070 70.445 146.135 ;
        RECT 70.735 146.120 70.965 146.210 ;
        RECT 68.530 145.840 70.530 146.070 ;
        RECT 68.610 145.775 70.445 145.840 ;
        RECT 71.725 145.100 72.725 152.410 ;
        RECT 74.900 146.775 75.900 157.100 ;
        RECT 85.530 152.775 86.530 153.310 ;
        RECT 88.600 153.295 89.600 157.100 ;
        RECT 77.125 152.450 78.980 152.570 ;
        RECT 82.410 152.450 84.260 152.575 ;
        RECT 77.050 152.220 79.050 152.450 ;
        RECT 82.335 152.220 84.335 152.450 ;
        RECT 85.480 152.410 86.530 152.775 ;
        RECT 77.125 152.210 78.980 152.220 ;
        RECT 82.410 152.215 84.260 152.220 ;
        RECT 76.660 151.840 76.890 152.170 ;
        RECT 79.210 151.840 79.440 152.170 ;
        RECT 80.185 151.840 81.145 151.870 ;
        RECT 81.900 151.840 82.130 152.170 ;
        RECT 84.540 151.840 84.770 152.170 ;
        RECT 76.660 151.540 84.770 151.840 ;
        RECT 76.660 151.210 76.890 151.540 ;
        RECT 79.210 151.210 79.440 151.540 ;
        RECT 80.185 151.510 81.145 151.540 ;
        RECT 81.900 151.210 82.130 151.540 ;
        RECT 84.540 151.210 84.770 151.540 ;
        RECT 77.050 150.930 79.050 151.160 ;
        RECT 82.335 150.930 84.335 151.160 ;
        RECT 77.105 150.790 78.995 150.930 ;
        RECT 82.390 150.790 84.280 150.930 ;
        RECT 77.105 150.590 84.280 150.790 ;
        RECT 77.125 150.020 78.975 150.150 ;
        RECT 77.050 149.790 79.050 150.020 ;
        RECT 76.660 149.650 76.890 149.740 ;
        RECT 79.210 149.650 79.440 149.740 ;
        RECT 80.755 149.650 81.155 150.590 ;
        RECT 82.410 150.020 84.255 150.155 ;
        RECT 82.335 149.790 84.335 150.020 ;
        RECT 81.900 149.650 82.130 149.740 ;
        RECT 84.540 149.650 84.770 149.740 ;
        RECT 76.660 149.440 84.770 149.650 ;
        RECT 76.660 149.370 76.980 149.440 ;
        RECT 79.120 149.370 82.270 149.440 ;
        RECT 84.405 149.370 84.770 149.440 ;
        RECT 76.660 149.280 76.890 149.370 ;
        RECT 77.125 149.230 78.975 149.295 ;
        RECT 79.210 149.280 79.440 149.370 ;
        RECT 77.050 149.000 79.050 149.230 ;
        RECT 76.660 148.860 76.890 148.950 ;
        RECT 77.125 148.935 78.975 149.000 ;
        RECT 79.210 148.860 79.440 148.950 ;
        RECT 80.755 148.860 81.155 149.370 ;
        RECT 81.900 149.280 82.130 149.370 ;
        RECT 82.415 149.230 84.260 149.295 ;
        RECT 84.540 149.280 84.770 149.370 ;
        RECT 82.335 149.000 84.335 149.230 ;
        RECT 81.900 148.860 82.130 148.950 ;
        RECT 82.415 148.935 84.260 149.000 ;
        RECT 84.540 148.860 84.770 148.950 ;
        RECT 76.660 148.790 76.980 148.860 ;
        RECT 79.120 148.790 82.270 148.860 ;
        RECT 84.405 148.790 84.770 148.860 ;
        RECT 76.660 148.650 84.770 148.790 ;
        RECT 76.660 148.580 76.980 148.650 ;
        RECT 79.120 148.580 82.270 148.650 ;
        RECT 84.405 148.580 84.770 148.650 ;
        RECT 76.660 148.490 76.890 148.580 ;
        RECT 77.130 148.440 78.975 148.505 ;
        RECT 79.210 148.490 79.440 148.580 ;
        RECT 77.050 148.210 79.050 148.440 ;
        RECT 76.660 148.070 76.890 148.160 ;
        RECT 77.130 148.145 78.975 148.210 ;
        RECT 79.210 148.070 79.440 148.160 ;
        RECT 80.755 148.070 81.155 148.580 ;
        RECT 81.900 148.490 82.130 148.580 ;
        RECT 82.425 148.440 84.275 148.505 ;
        RECT 84.540 148.490 84.770 148.580 ;
        RECT 82.335 148.210 84.335 148.440 ;
        RECT 81.900 148.070 82.130 148.160 ;
        RECT 82.425 148.145 84.275 148.210 ;
        RECT 84.540 148.070 84.770 148.160 ;
        RECT 76.660 148.000 76.980 148.070 ;
        RECT 79.120 148.000 82.270 148.070 ;
        RECT 84.405 148.000 84.770 148.070 ;
        RECT 76.660 147.860 84.770 148.000 ;
        RECT 76.660 147.790 76.985 147.860 ;
        RECT 79.120 147.790 82.270 147.860 ;
        RECT 84.405 147.790 84.770 147.860 ;
        RECT 76.660 147.700 76.890 147.790 ;
        RECT 77.130 147.650 78.975 147.715 ;
        RECT 79.210 147.700 79.440 147.790 ;
        RECT 77.050 147.420 79.050 147.650 ;
        RECT 77.130 147.355 78.975 147.420 ;
        RECT 81.435 147.280 81.695 147.790 ;
        RECT 81.900 147.700 82.130 147.790 ;
        RECT 82.425 147.650 84.250 147.715 ;
        RECT 84.540 147.700 84.770 147.790 ;
        RECT 82.335 147.420 84.335 147.650 ;
        RECT 81.900 147.280 82.130 147.370 ;
        RECT 82.425 147.355 84.250 147.420 ;
        RECT 84.540 147.280 84.770 147.370 ;
        RECT 81.435 147.210 82.270 147.280 ;
        RECT 84.405 147.210 84.770 147.280 ;
        RECT 81.435 147.070 84.770 147.210 ;
        RECT 81.435 147.000 82.270 147.070 ;
        RECT 84.405 147.000 84.770 147.070 ;
        RECT 81.435 146.490 81.695 147.000 ;
        RECT 81.900 146.910 82.130 147.000 ;
        RECT 82.410 146.860 84.260 146.925 ;
        RECT 84.540 146.910 84.770 147.000 ;
        RECT 82.335 146.630 84.335 146.860 ;
        RECT 81.900 146.490 82.130 146.580 ;
        RECT 82.410 146.565 84.260 146.630 ;
        RECT 84.540 146.490 84.770 146.580 ;
        RECT 81.435 146.420 82.270 146.490 ;
        RECT 84.405 146.420 84.770 146.490 ;
        RECT 81.435 146.280 84.770 146.420 ;
        RECT 81.435 146.210 82.270 146.280 ;
        RECT 84.405 146.210 84.770 146.280 ;
        RECT 81.900 146.120 82.130 146.210 ;
        RECT 82.415 146.070 84.250 146.135 ;
        RECT 84.540 146.120 84.770 146.210 ;
        RECT 82.335 145.840 84.335 146.070 ;
        RECT 82.415 145.775 84.250 145.840 ;
        RECT 85.530 145.100 86.530 152.410 ;
        RECT 88.590 153.100 89.600 153.295 ;
        RECT 88.590 146.775 89.590 153.100 ;
        RECT 99.220 152.775 100.220 153.310 ;
        RECT 90.815 152.450 92.670 152.570 ;
        RECT 96.100 152.450 97.950 152.575 ;
        RECT 90.740 152.220 92.740 152.450 ;
        RECT 96.025 152.220 98.025 152.450 ;
        RECT 99.170 152.410 100.220 152.775 ;
        RECT 90.815 152.210 92.670 152.220 ;
        RECT 96.100 152.215 97.950 152.220 ;
        RECT 90.350 151.840 90.580 152.170 ;
        RECT 92.900 151.840 93.130 152.170 ;
        RECT 93.875 151.840 94.835 151.870 ;
        RECT 95.590 151.840 95.820 152.170 ;
        RECT 98.230 151.840 98.460 152.170 ;
        RECT 90.350 151.540 98.460 151.840 ;
        RECT 90.350 151.210 90.580 151.540 ;
        RECT 92.900 151.210 93.130 151.540 ;
        RECT 93.875 151.510 94.835 151.540 ;
        RECT 95.590 151.210 95.820 151.540 ;
        RECT 98.230 151.210 98.460 151.540 ;
        RECT 90.740 150.930 92.740 151.160 ;
        RECT 96.025 150.930 98.025 151.160 ;
        RECT 90.795 150.790 92.685 150.930 ;
        RECT 96.080 150.790 97.970 150.930 ;
        RECT 90.795 150.590 97.970 150.790 ;
        RECT 90.815 150.020 92.665 150.150 ;
        RECT 90.740 149.790 92.740 150.020 ;
        RECT 90.350 149.650 90.580 149.740 ;
        RECT 92.900 149.650 93.130 149.740 ;
        RECT 94.445 149.650 94.845 150.590 ;
        RECT 96.100 150.020 97.945 150.155 ;
        RECT 96.025 149.790 98.025 150.020 ;
        RECT 95.590 149.650 95.820 149.740 ;
        RECT 98.230 149.650 98.460 149.740 ;
        RECT 90.350 149.440 98.460 149.650 ;
        RECT 90.350 149.370 90.670 149.440 ;
        RECT 92.810 149.370 95.960 149.440 ;
        RECT 98.095 149.370 98.460 149.440 ;
        RECT 90.350 149.280 90.580 149.370 ;
        RECT 90.815 149.230 92.665 149.295 ;
        RECT 92.900 149.280 93.130 149.370 ;
        RECT 90.740 149.000 92.740 149.230 ;
        RECT 90.350 148.860 90.580 148.950 ;
        RECT 90.815 148.935 92.665 149.000 ;
        RECT 92.900 148.860 93.130 148.950 ;
        RECT 94.445 148.860 94.845 149.370 ;
        RECT 95.590 149.280 95.820 149.370 ;
        RECT 96.105 149.230 97.950 149.295 ;
        RECT 98.230 149.280 98.460 149.370 ;
        RECT 96.025 149.000 98.025 149.230 ;
        RECT 95.590 148.860 95.820 148.950 ;
        RECT 96.105 148.935 97.950 149.000 ;
        RECT 98.230 148.860 98.460 148.950 ;
        RECT 90.350 148.790 90.670 148.860 ;
        RECT 92.810 148.790 95.960 148.860 ;
        RECT 98.095 148.790 98.460 148.860 ;
        RECT 90.350 148.650 98.460 148.790 ;
        RECT 90.350 148.580 90.670 148.650 ;
        RECT 92.810 148.580 95.960 148.650 ;
        RECT 98.095 148.580 98.460 148.650 ;
        RECT 90.350 148.490 90.580 148.580 ;
        RECT 90.820 148.440 92.665 148.505 ;
        RECT 92.900 148.490 93.130 148.580 ;
        RECT 90.740 148.210 92.740 148.440 ;
        RECT 90.350 148.070 90.580 148.160 ;
        RECT 90.820 148.145 92.665 148.210 ;
        RECT 92.900 148.070 93.130 148.160 ;
        RECT 94.445 148.070 94.845 148.580 ;
        RECT 95.590 148.490 95.820 148.580 ;
        RECT 96.115 148.440 97.965 148.505 ;
        RECT 98.230 148.490 98.460 148.580 ;
        RECT 96.025 148.210 98.025 148.440 ;
        RECT 95.590 148.070 95.820 148.160 ;
        RECT 96.115 148.145 97.965 148.210 ;
        RECT 98.230 148.070 98.460 148.160 ;
        RECT 90.350 148.000 90.670 148.070 ;
        RECT 92.810 148.000 95.960 148.070 ;
        RECT 98.095 148.000 98.460 148.070 ;
        RECT 90.350 147.860 98.460 148.000 ;
        RECT 90.350 147.790 90.675 147.860 ;
        RECT 92.810 147.790 95.960 147.860 ;
        RECT 98.095 147.790 98.460 147.860 ;
        RECT 90.350 147.700 90.580 147.790 ;
        RECT 90.820 147.650 92.665 147.715 ;
        RECT 92.900 147.700 93.130 147.790 ;
        RECT 90.740 147.420 92.740 147.650 ;
        RECT 90.820 147.355 92.665 147.420 ;
        RECT 95.125 147.280 95.385 147.790 ;
        RECT 95.590 147.700 95.820 147.790 ;
        RECT 96.115 147.650 97.940 147.715 ;
        RECT 98.230 147.700 98.460 147.790 ;
        RECT 96.025 147.420 98.025 147.650 ;
        RECT 95.590 147.280 95.820 147.370 ;
        RECT 96.115 147.355 97.940 147.420 ;
        RECT 98.230 147.280 98.460 147.370 ;
        RECT 95.125 147.210 95.960 147.280 ;
        RECT 98.095 147.210 98.460 147.280 ;
        RECT 95.125 147.070 98.460 147.210 ;
        RECT 95.125 147.000 95.960 147.070 ;
        RECT 98.095 147.000 98.460 147.070 ;
        RECT 95.125 146.490 95.385 147.000 ;
        RECT 95.590 146.910 95.820 147.000 ;
        RECT 96.100 146.860 97.950 146.925 ;
        RECT 98.230 146.910 98.460 147.000 ;
        RECT 96.025 146.630 98.025 146.860 ;
        RECT 95.590 146.490 95.820 146.580 ;
        RECT 96.100 146.565 97.950 146.630 ;
        RECT 98.230 146.490 98.460 146.580 ;
        RECT 95.125 146.420 95.960 146.490 ;
        RECT 98.095 146.420 98.460 146.490 ;
        RECT 95.125 146.280 98.460 146.420 ;
        RECT 95.125 146.210 95.960 146.280 ;
        RECT 98.095 146.210 98.460 146.280 ;
        RECT 95.590 146.120 95.820 146.210 ;
        RECT 96.105 146.070 97.940 146.135 ;
        RECT 98.230 146.120 98.460 146.210 ;
        RECT 96.025 145.840 98.025 146.070 ;
        RECT 96.105 145.775 97.940 145.840 ;
        RECT 99.220 145.100 100.220 152.410 ;
        RECT 58.195 145.060 59.200 145.100 ;
        RECT 58.200 141.500 59.200 145.060 ;
        RECT 71.700 145.035 72.725 145.100 ;
        RECT 85.500 145.035 86.530 145.100 ;
        RECT 99.200 145.035 100.220 145.100 ;
        RECT 71.700 141.500 72.700 145.035 ;
        RECT 67.285 135.950 67.535 138.055 ;
        RECT 69.290 136.190 69.540 136.255 ;
        RECT 69.235 134.240 69.595 136.190 ;
        RECT 75.320 135.990 75.570 136.055 ;
        RECT 71.300 135.790 71.550 135.855 ;
        RECT 73.310 135.790 73.560 135.855 ;
        RECT 69.290 134.150 69.540 134.240 ;
        RECT 71.245 133.840 71.605 135.790 ;
        RECT 73.255 133.840 73.615 135.790 ;
        RECT 75.265 134.040 75.625 135.990 ;
        RECT 75.320 133.950 75.570 134.040 ;
        RECT 71.300 133.750 71.550 133.840 ;
        RECT 73.310 133.750 73.560 133.840 ;
        RECT 67.285 123.985 67.535 124.060 ;
        RECT 69.290 123.985 69.540 124.060 ;
        RECT 71.300 123.995 71.550 124.060 ;
        RECT 73.310 123.995 73.560 124.060 ;
        RECT 75.320 123.995 75.570 124.060 ;
        RECT 67.240 122.035 67.600 123.985 ;
        RECT 69.190 122.035 69.550 123.985 ;
        RECT 71.245 122.045 71.605 123.995 ;
        RECT 73.255 122.045 73.615 123.995 ;
        RECT 75.265 122.045 75.625 123.995 ;
        RECT 82.300 122.500 83.300 144.000 ;
        RECT 85.500 141.500 86.500 145.035 ;
        RECT 99.200 141.500 100.200 145.035 ;
        RECT 104.600 137.690 105.600 156.400 ;
        RECT 85.320 136.475 114.300 137.690 ;
        RECT 85.810 136.400 86.990 136.475 ;
        RECT 88.085 135.805 92.045 136.035 ;
        RECT 87.805 133.555 88.035 135.645 ;
        RECT 87.620 132.440 88.035 133.555 ;
        RECT 87.805 131.645 88.035 132.440 ;
        RECT 89.300 131.485 90.820 135.805 ;
        RECT 92.400 135.650 93.185 136.475 ;
        RECT 93.515 135.805 97.475 136.035 ;
        RECT 101.125 136.000 102.985 136.475 ;
        RECT 104.690 136.000 106.535 136.475 ;
        RECT 92.145 135.645 93.420 135.650 ;
        RECT 92.095 134.375 93.465 135.645 ;
        RECT 92.095 131.645 92.325 134.375 ;
        RECT 93.235 131.645 93.465 134.375 ;
        RECT 94.820 134.550 96.340 135.805 ;
        RECT 101.045 135.770 103.045 136.000 ;
        RECT 104.615 135.770 106.615 136.000 ;
        RECT 97.525 134.550 97.755 135.645 ;
        RECT 94.820 134.490 97.755 134.550 ;
        RECT 94.820 132.955 99.545 134.490 ;
        RECT 100.655 134.260 100.885 135.720 ;
        RECT 100.500 134.190 100.885 134.260 ;
        RECT 103.205 134.190 103.435 135.720 ;
        RECT 100.500 133.195 103.435 134.190 ;
        RECT 94.820 132.935 97.755 132.955 ;
        RECT 94.820 131.485 96.340 132.935 ;
        RECT 97.525 131.645 97.755 132.935 ;
        RECT 88.085 131.255 92.045 131.485 ;
        RECT 93.515 131.255 97.475 131.485 ;
        RECT 98.520 129.455 99.525 132.955 ;
        RECT 100.500 132.945 100.885 133.195 ;
        RECT 100.655 131.760 100.885 132.945 ;
        RECT 103.205 131.760 103.435 133.195 ;
        RECT 104.225 134.185 104.455 135.720 ;
        RECT 106.775 134.185 107.005 135.720 ;
        RECT 104.225 133.205 108.945 134.185 ;
        RECT 109.140 133.585 109.895 136.475 ;
        RECT 110.905 133.820 111.365 134.050 ;
        RECT 110.985 133.800 111.240 133.820 ;
        RECT 110.625 133.585 110.855 133.660 ;
        RECT 104.225 133.185 107.005 133.205 ;
        RECT 104.225 131.760 104.455 133.185 ;
        RECT 106.775 131.760 107.005 133.185 ;
        RECT 101.045 131.480 103.045 131.710 ;
        RECT 104.615 131.480 106.615 131.710 ;
        RECT 101.075 131.355 103.015 131.480 ;
        RECT 104.650 131.355 106.605 131.480 ;
        RECT 107.805 129.455 108.945 133.205 ;
        RECT 109.125 133.110 110.855 133.585 ;
        RECT 110.625 133.050 110.855 133.110 ;
        RECT 111.010 132.905 111.240 133.800 ;
        RECT 111.415 133.600 111.645 133.660 ;
        RECT 111.415 133.135 113.905 133.600 ;
        RECT 111.415 133.050 111.645 133.135 ;
        RECT 110.985 132.890 111.240 132.905 ;
        RECT 110.905 132.660 111.365 132.890 ;
        RECT 110.980 129.725 111.240 132.660 ;
        RECT 98.520 129.450 108.945 129.455 ;
        RECT 94.520 129.395 108.945 129.450 ;
        RECT 94.495 128.590 108.945 129.395 ;
        RECT 109.940 128.785 111.240 129.725 ;
        RECT 88.090 127.300 90.050 127.530 ;
        RECT 91.520 127.300 93.480 127.530 ;
        RECT 87.810 126.850 88.040 127.095 ;
        RECT 87.670 125.690 88.050 126.850 ;
        RECT 87.810 123.095 88.040 125.690 ;
        RECT 88.785 122.965 89.445 127.300 ;
        RECT 90.100 125.880 90.330 127.095 ;
        RECT 91.240 125.880 91.470 127.095 ;
        RECT 90.100 123.095 91.470 125.880 ;
        RECT 88.115 122.890 90.020 122.965 ;
        RECT 88.090 122.660 90.050 122.890 ;
        RECT 82.300 122.320 85.900 122.500 ;
        RECT 82.300 122.285 86.790 122.320 ;
        RECT 90.190 122.285 91.320 123.095 ;
        RECT 92.155 122.955 92.815 127.300 ;
        RECT 93.530 125.630 93.760 127.095 ;
        RECT 94.495 125.630 95.805 128.590 ;
        RECT 97.135 127.295 99.095 127.525 ;
        RECT 99.425 127.295 101.385 127.525 ;
        RECT 102.855 127.295 104.815 127.525 ;
        RECT 105.145 127.295 107.105 127.525 ;
        RECT 93.530 124.140 95.810 125.630 ;
        RECT 96.855 125.470 97.085 127.090 ;
        RECT 96.830 124.580 97.200 125.470 ;
        RECT 93.530 123.095 93.760 124.140 ;
        RECT 96.855 123.090 97.085 124.580 ;
        RECT 91.565 122.890 93.470 122.955 ;
        RECT 91.520 122.660 93.480 122.890 ;
        RECT 97.670 122.885 98.650 127.295 ;
        RECT 99.145 126.975 99.375 127.090 ;
        RECT 99.125 125.855 99.490 126.975 ;
        RECT 99.145 123.090 99.375 125.855 ;
        RECT 99.995 122.885 100.935 127.295 ;
        RECT 101.435 125.475 101.665 127.090 ;
        RECT 102.575 125.505 102.805 127.090 ;
        RECT 101.270 124.570 101.680 125.475 ;
        RECT 102.550 124.585 102.920 125.505 ;
        RECT 101.435 123.090 101.665 124.570 ;
        RECT 102.575 123.090 102.805 124.585 ;
        RECT 103.330 122.885 104.285 127.295 ;
        RECT 104.865 126.995 105.095 127.090 ;
        RECT 104.845 125.935 105.240 126.995 ;
        RECT 104.865 123.090 105.095 125.935 ;
        RECT 105.635 122.885 106.590 127.295 ;
        RECT 107.155 125.505 107.385 127.090 ;
        RECT 110.980 126.520 111.240 128.785 ;
        RECT 110.880 126.290 111.340 126.520 ;
        RECT 114.800 126.400 125.300 127.400 ;
        RECT 110.600 126.030 110.830 126.085 ;
        RECT 107.020 124.580 107.385 125.505 ;
        RECT 107.155 123.090 107.385 124.580 ;
        RECT 109.000 125.640 110.830 126.030 ;
        RECT 97.135 122.655 99.095 122.885 ;
        RECT 99.425 122.655 101.385 122.885 ;
        RECT 102.855 122.655 104.815 122.885 ;
        RECT 105.145 122.655 107.105 122.885 ;
        RECT 109.000 122.285 109.695 125.640 ;
        RECT 110.600 125.585 110.830 125.640 ;
        RECT 110.980 125.380 111.220 126.290 ;
        RECT 111.390 126.040 111.620 126.085 ;
        RECT 111.390 125.650 113.920 126.040 ;
        RECT 111.390 125.585 111.620 125.650 ;
        RECT 110.880 125.150 111.340 125.380 ;
        RECT 114.800 125.100 115.800 126.400 ;
        RECT 113.200 124.100 115.800 125.100 ;
        RECT 124.300 125.000 125.300 126.400 ;
        RECT 113.200 122.285 114.300 124.100 ;
        RECT 120.355 124.090 121.315 124.320 ;
        RECT 67.285 121.955 67.535 122.035 ;
        RECT 69.290 121.955 69.540 122.035 ;
        RECT 71.300 121.955 71.550 122.045 ;
        RECT 73.310 121.955 73.560 122.045 ;
        RECT 75.320 121.955 75.570 122.045 ;
        RECT 82.300 120.900 114.300 122.285 ;
        RECT 120.075 121.875 120.305 123.885 ;
        RECT 85.300 120.860 114.300 120.900 ;
        RECT 66.830 111.020 67.830 120.555 ;
        RECT 69.290 120.170 69.540 120.235 ;
        RECT 71.300 120.170 71.550 120.235 ;
        RECT 73.310 120.170 73.560 120.235 ;
        RECT 69.235 118.220 69.595 120.170 ;
        RECT 71.245 118.220 71.605 120.170 ;
        RECT 73.255 118.220 73.615 120.170 ;
        RECT 119.970 119.950 120.330 121.875 ;
        RECT 120.075 119.885 120.305 119.950 ;
        RECT 120.680 119.680 120.980 124.090 ;
        RECT 122.415 124.000 125.295 125.000 ;
        RECT 121.365 121.860 121.595 123.885 ;
        RECT 122.615 122.010 123.070 122.610 ;
        RECT 121.345 119.940 121.745 121.860 ;
        RECT 123.315 121.090 124.275 121.320 ;
        RECT 123.035 120.810 123.265 120.885 ;
        RECT 122.915 119.955 123.275 120.810 ;
        RECT 121.365 119.885 121.595 119.940 ;
        RECT 123.035 119.885 123.265 119.955 ;
        RECT 123.640 119.680 123.940 121.090 ;
        RECT 124.325 120.810 124.555 120.885 ;
        RECT 124.310 119.950 124.680 120.810 ;
        RECT 124.325 119.885 124.555 119.950 ;
        RECT 120.355 119.450 121.315 119.680 ;
        RECT 123.315 119.450 124.275 119.680 ;
        RECT 120.680 118.575 120.980 119.450 ;
        RECT 120.675 118.245 120.980 118.575 ;
        RECT 123.640 118.320 123.940 119.450 ;
        RECT 122.885 118.295 123.940 118.320 ;
        RECT 120.585 118.225 120.980 118.245 ;
        RECT 69.290 118.130 69.540 118.220 ;
        RECT 71.300 118.130 71.550 118.220 ;
        RECT 73.310 118.130 73.560 118.220 ;
        RECT 120.565 117.965 120.980 118.225 ;
        RECT 120.585 117.945 120.980 117.965 ;
        RECT 122.865 117.950 123.940 118.295 ;
        RECT 120.675 117.615 120.980 117.945 ;
        RECT 122.885 117.920 123.940 117.950 ;
        RECT 120.680 116.820 120.980 117.615 ;
        RECT 123.640 116.820 123.940 117.920 ;
        RECT 120.350 116.590 121.310 116.820 ;
        RECT 123.310 116.590 124.270 116.820 ;
        RECT 120.070 116.370 120.300 116.430 ;
        RECT 77.000 115.660 82.100 115.700 ;
        RECT 77.000 114.660 101.855 115.660 ;
        RECT 77.000 114.600 82.100 114.660 ;
        RECT 69.290 113.375 69.540 113.440 ;
        RECT 71.300 113.375 71.550 113.440 ;
        RECT 73.310 113.375 73.560 113.440 ;
        RECT 69.235 111.425 69.595 113.375 ;
        RECT 71.245 111.425 71.605 113.375 ;
        RECT 73.255 111.425 73.615 113.375 ;
        RECT 69.290 111.335 69.540 111.425 ;
        RECT 71.300 111.335 71.550 111.425 ;
        RECT 73.310 111.335 73.560 111.425 ;
        RECT 77.000 109.000 78.200 114.600 ;
        RECT 83.220 113.610 85.180 113.840 ;
        RECT 90.170 113.610 91.130 113.840 ;
        RECT 82.940 113.320 83.170 113.405 ;
        RECT 82.875 111.410 83.235 113.320 ;
        RECT 82.940 109.405 83.170 111.410 ;
        RECT 84.055 109.200 84.355 113.610 ;
        RECT 85.230 109.405 85.460 113.405 ;
        RECT 89.890 111.390 90.120 113.405 ;
        RECT 89.755 109.485 90.120 111.390 ;
        RECT 89.890 109.405 90.120 109.485 ;
        RECT 90.500 109.200 90.800 113.610 ;
        RECT 91.180 113.355 91.410 113.405 ;
        RECT 91.615 113.355 92.115 114.660 ;
        RECT 119.970 114.475 120.330 116.370 ;
        RECT 92.600 113.610 93.560 113.840 ;
        RECT 98.560 113.615 100.520 113.845 ;
        RECT 92.320 113.355 92.550 113.405 ;
        RECT 91.180 111.385 92.550 113.355 ;
        RECT 91.180 109.405 91.410 111.385 ;
        RECT 92.320 109.405 92.550 111.385 ;
        RECT 92.930 109.200 93.230 113.610 ;
        RECT 93.610 111.405 93.840 113.405 ;
        RECT 93.610 109.490 93.975 111.405 ;
        RECT 93.610 109.405 93.840 109.490 ;
        RECT 98.280 109.410 98.510 113.410 ;
        RECT 99.390 109.205 99.690 113.615 ;
        RECT 100.570 113.330 100.800 113.410 ;
        RECT 100.505 111.415 100.865 113.330 ;
        RECT 120.070 112.430 120.300 114.475 ;
        RECT 120.680 112.270 120.980 116.590 ;
        RECT 121.360 116.365 121.590 116.430 ;
        RECT 121.350 114.445 121.750 116.365 ;
        RECT 123.030 116.355 123.260 116.430 ;
        RECT 122.910 115.495 123.270 116.355 ;
        RECT 123.030 115.430 123.260 115.495 ;
        RECT 123.640 115.270 123.940 116.590 ;
        RECT 124.320 116.345 124.550 116.430 ;
        RECT 124.315 115.515 124.685 116.345 ;
        RECT 124.320 115.430 124.550 115.515 ;
        RECT 123.310 115.040 124.270 115.270 ;
        RECT 121.360 112.430 121.590 114.445 ;
        RECT 122.620 113.880 123.080 114.495 ;
        RECT 120.350 112.040 121.310 112.270 ;
        RECT 100.570 109.410 100.800 111.415 ;
        RECT 122.460 111.400 125.265 112.320 ;
        RECT 122.460 111.320 125.300 111.400 ;
        RECT 104.810 110.630 105.270 110.860 ;
        RECT 104.530 109.925 104.760 110.425 ;
        RECT 104.910 109.720 105.170 110.630 ;
        RECT 105.320 110.360 105.550 110.425 ;
        RECT 105.320 109.990 105.680 110.360 ;
        RECT 105.320 109.925 105.550 109.990 ;
        RECT 104.810 109.490 105.270 109.720 ;
        RECT 46.500 108.000 78.200 109.000 ;
        RECT 83.220 108.970 85.180 109.200 ;
        RECT 90.170 108.970 91.130 109.200 ;
        RECT 92.600 108.970 93.560 109.200 ;
        RECT 98.560 108.975 100.520 109.205 ;
        RECT 84.830 108.190 85.130 108.970 ;
        RECT 90.230 108.190 90.580 108.970 ;
        RECT 93.145 108.195 93.505 108.970 ;
        RECT 98.615 108.195 98.915 108.975 ;
        RECT 84.795 107.930 85.165 108.190 ;
        RECT 90.195 107.930 90.610 108.190 ;
        RECT 93.110 107.935 93.540 108.195 ;
        RECT 98.580 107.935 98.950 108.195 ;
        RECT 104.910 108.145 105.170 109.490 ;
        RECT 100.505 107.885 105.170 108.145 ;
        RECT 82.875 107.500 98.915 107.760 ;
        RECT 82.830 106.990 83.280 107.005 ;
        RECT 80.930 106.760 85.180 106.990 ;
        RECT 98.615 106.985 98.915 107.500 ;
        RECT 104.910 106.985 105.170 107.885 ;
        RECT 98.560 106.960 100.520 106.985 ;
        RECT 100.850 106.960 102.810 106.985 ;
        RECT 98.560 106.780 102.810 106.960 ;
        RECT 80.650 102.600 80.880 106.600 ;
        RECT 81.760 102.440 82.060 106.760 ;
        RECT 82.830 106.745 83.280 106.760 ;
        RECT 82.940 104.605 83.170 106.600 ;
        RECT 82.875 102.695 83.235 104.605 ;
        RECT 82.940 102.600 83.170 102.695 ;
        RECT 84.050 102.440 84.350 106.760 ;
        RECT 98.560 106.755 100.520 106.780 ;
        RECT 100.850 106.755 102.810 106.780 ;
        RECT 104.810 106.755 105.270 106.985 ;
        RECT 85.230 102.600 85.460 106.600 ;
        RECT 89.005 106.410 89.505 106.465 ;
        RECT 94.020 106.415 94.520 106.475 ;
        RECT 88.985 106.110 89.525 106.410 ;
        RECT 94.010 106.115 94.525 106.415 ;
        RECT 89.005 104.990 89.505 106.110 ;
        RECT 94.020 104.990 94.520 106.115 ;
        RECT 87.170 104.760 91.130 104.990 ;
        RECT 92.600 104.760 96.560 104.990 ;
        RECT 86.890 104.520 87.120 104.600 ;
        RECT 86.755 102.690 87.120 104.520 ;
        RECT 86.890 102.600 87.120 102.690 ;
        RECT 89.005 102.440 89.505 104.760 ;
        RECT 91.180 104.545 91.410 104.600 ;
        RECT 92.320 104.545 92.550 104.600 ;
        RECT 91.180 102.655 92.550 104.545 ;
        RECT 91.180 102.600 91.410 102.655 ;
        RECT 80.930 102.415 82.890 102.440 ;
        RECT 83.220 102.415 85.180 102.440 ;
        RECT 80.930 102.210 85.180 102.415 ;
        RECT 87.170 102.210 91.130 102.440 ;
        RECT 91.615 101.205 92.115 102.655 ;
        RECT 92.320 102.600 92.550 102.655 ;
        RECT 94.020 102.440 94.520 104.760 ;
        RECT 96.610 104.520 96.840 104.600 ;
        RECT 96.610 102.685 96.975 104.520 ;
        RECT 96.610 102.600 96.840 102.685 ;
        RECT 98.280 102.595 98.510 106.595 ;
        RECT 92.600 102.210 96.560 102.440 ;
        RECT 99.390 102.435 99.690 106.755 ;
        RECT 100.570 104.595 100.800 106.595 ;
        RECT 100.505 102.680 100.865 104.595 ;
        RECT 100.570 102.595 100.800 102.680 ;
        RECT 101.680 102.435 101.980 106.755 ;
        RECT 102.860 102.595 103.090 106.595 ;
        RECT 104.530 104.795 104.760 106.595 ;
        RECT 104.910 104.635 105.170 106.755 ;
        RECT 105.320 106.525 105.550 106.595 ;
        RECT 105.320 105.705 105.690 106.525 ;
        RECT 105.320 104.795 105.550 105.705 ;
        RECT 104.810 104.405 105.270 104.635 ;
        RECT 98.560 102.410 100.520 102.435 ;
        RECT 100.850 102.410 102.810 102.435 ;
        RECT 98.560 102.230 102.810 102.410 ;
        RECT 98.560 102.205 100.520 102.230 ;
        RECT 100.850 102.205 102.810 102.230 ;
        RECT 79.850 101.200 105.530 101.205 ;
        RECT 124.300 101.200 125.300 111.320 ;
        RECT 79.850 100.205 125.300 101.200 ;
        RECT 105.400 100.200 125.300 100.205 ;
      LAYER met2 ;
        RECT 72.700 184.500 73.300 219.200 ;
        RECT 77.700 217.300 78.900 217.900 ;
        RECT 140.800 213.600 141.500 213.700 ;
        RECT 105.200 213.000 141.500 213.600 ;
        RECT 105.200 211.000 105.800 213.000 ;
        RECT 143.600 211.000 144.300 211.100 ;
        RECT 94.900 210.400 105.800 211.000 ;
        RECT 115.200 210.500 144.300 211.000 ;
        RECT 95.080 207.410 95.360 210.400 ;
        RECT 115.320 207.410 115.600 210.500 ;
        RECT 143.600 210.400 144.300 210.500 ;
        RECT 95.080 207.270 95.750 207.410 ;
        RECT 95.080 206.755 95.360 207.270 ;
        RECT 92.320 203.075 92.600 203.445 ;
        RECT 92.390 197.130 92.530 203.075 ;
        RECT 92.330 196.810 92.590 197.130 ;
        RECT 95.610 196.450 95.750 207.270 ;
        RECT 115.320 207.270 115.990 207.410 ;
        RECT 115.320 206.755 115.600 207.270 ;
        RECT 98.610 197.295 100.490 197.665 ;
        RECT 106.110 197.295 107.990 197.665 ;
        RECT 113.610 197.295 115.490 197.665 ;
        RECT 95.550 196.130 95.810 196.450 ;
        RECT 101.070 195.790 101.330 196.110 ;
        RECT 93.710 195.110 93.970 195.430 ;
        RECT 100.610 195.110 100.870 195.430 ;
        RECT 93.770 193.925 93.910 195.110 ;
        RECT 94.910 194.575 96.790 194.945 ;
        RECT 93.700 193.555 93.980 193.925 ;
        RECT 98.610 191.855 100.490 192.225 ;
        RECT 99.690 190.350 99.950 190.670 ;
        RECT 94.910 189.135 96.790 189.505 ;
        RECT 93.250 187.630 93.510 187.950 ;
        RECT 89.560 184.715 89.840 185.085 ;
        RECT 89.630 184.550 89.770 184.715 ;
        RECT 89.570 184.230 89.830 184.550 ;
        RECT 93.310 182.510 93.450 187.630 ;
        RECT 99.750 187.270 99.890 190.350 ;
        RECT 100.670 188.970 100.810 195.110 ;
        RECT 100.610 188.650 100.870 188.970 ;
        RECT 100.610 187.970 100.870 188.290 ;
        RECT 99.690 186.950 99.950 187.270 ;
        RECT 98.610 186.415 100.490 186.785 ;
        RECT 97.390 185.250 97.650 185.570 ;
        RECT 94.910 183.695 96.790 184.065 ;
        RECT 97.450 183.530 97.590 185.250 ;
        RECT 97.390 183.210 97.650 183.530 ;
        RECT 93.250 182.190 93.510 182.510 ;
        RECT 93.310 177.070 93.450 182.190 ;
        RECT 97.450 180.810 97.590 183.210 ;
        RECT 97.850 181.850 98.110 182.170 ;
        RECT 97.390 180.490 97.650 180.810 ;
        RECT 97.910 180.130 98.050 181.850 ;
        RECT 98.610 180.975 100.490 181.345 ;
        RECT 97.850 179.810 98.110 180.130 ;
        RECT 94.910 178.255 96.790 178.625 ;
        RECT 100.670 177.750 100.810 187.970 ;
        RECT 101.130 186.250 101.270 195.790 ;
        RECT 105.670 195.450 105.930 195.770 ;
        RECT 102.410 194.575 104.290 194.945 ;
        RECT 104.750 191.030 105.010 191.350 ;
        RECT 102.410 189.135 104.290 189.505 ;
        RECT 104.810 188.970 104.950 191.030 ;
        RECT 105.210 190.010 105.470 190.330 ;
        RECT 104.750 188.650 105.010 188.970 ;
        RECT 105.270 188.370 105.410 190.010 ;
        RECT 105.730 188.970 105.870 195.450 ;
        RECT 109.910 194.575 111.790 194.945 ;
        RECT 108.890 192.730 109.150 193.050 ;
        RECT 106.110 191.855 107.990 192.225 ;
        RECT 105.670 188.650 105.930 188.970 ;
        RECT 105.270 188.230 105.870 188.370 ;
        RECT 105.730 187.610 105.870 188.230 ;
        RECT 101.990 187.290 102.250 187.610 ;
        RECT 105.210 187.290 105.470 187.610 ;
        RECT 105.670 187.290 105.930 187.610 ;
        RECT 101.070 185.930 101.330 186.250 ;
        RECT 101.130 182.930 101.270 185.930 ;
        RECT 102.050 185.570 102.190 187.290 ;
        RECT 104.750 186.950 105.010 187.270 ;
        RECT 101.990 185.250 102.250 185.570 ;
        RECT 104.810 184.970 104.950 186.950 ;
        RECT 105.270 185.910 105.410 187.290 ;
        RECT 105.210 185.590 105.470 185.910 ;
        RECT 104.810 184.830 105.410 184.970 ;
        RECT 105.730 184.890 105.870 187.290 ;
        RECT 106.110 186.415 107.990 186.785 ;
        RECT 108.430 184.910 108.690 185.230 ;
        RECT 102.410 183.695 104.290 184.065 ;
        RECT 101.130 182.790 101.730 182.930 ;
        RECT 101.070 182.190 101.330 182.510 ;
        RECT 100.610 177.430 100.870 177.750 ;
        RECT 101.130 177.410 101.270 182.190 ;
        RECT 101.590 180.810 101.730 182.790 ;
        RECT 104.750 182.530 105.010 182.850 ;
        RECT 104.290 182.190 104.550 182.510 ;
        RECT 101.530 180.490 101.790 180.810 ;
        RECT 101.990 180.150 102.250 180.470 ;
        RECT 101.530 179.810 101.790 180.130 ;
        RECT 101.590 179.110 101.730 179.810 ;
        RECT 101.530 178.790 101.790 179.110 ;
        RECT 101.070 177.090 101.330 177.410 ;
        RECT 93.250 176.750 93.510 177.070 ;
        RECT 77.700 174.400 78.300 176.600 ;
        RECT 89.560 173.835 89.840 174.205 ;
        RECT 89.570 173.690 89.830 173.835 ;
        RECT 93.310 172.650 93.450 176.750 ;
        RECT 101.590 176.730 101.730 178.790 ;
        RECT 102.050 177.070 102.190 180.150 ;
        RECT 104.350 179.110 104.490 182.190 ;
        RECT 104.290 178.790 104.550 179.110 ;
        RECT 102.410 178.255 104.290 178.625 ;
        RECT 104.810 178.090 104.950 182.530 ;
        RECT 104.750 177.770 105.010 178.090 ;
        RECT 105.270 177.490 105.410 184.830 ;
        RECT 105.670 184.570 105.930 184.890 ;
        RECT 105.730 182.510 105.870 184.570 ;
        RECT 105.670 182.190 105.930 182.510 ;
        RECT 105.670 181.510 105.930 181.830 ;
        RECT 104.810 177.410 105.410 177.490 ;
        RECT 104.750 177.350 105.410 177.410 ;
        RECT 104.750 177.090 105.010 177.350 ;
        RECT 101.990 176.750 102.250 177.070 ;
        RECT 101.530 176.410 101.790 176.730 ;
        RECT 98.610 175.535 100.490 175.905 ;
        RECT 101.590 174.770 101.730 176.410 ;
        RECT 101.130 174.690 101.730 174.770 ;
        RECT 101.070 174.630 101.730 174.690 ;
        RECT 101.070 174.370 101.330 174.630 ;
        RECT 93.710 173.350 93.970 173.670 ;
        RECT 93.250 172.330 93.510 172.650 ;
        RECT 93.770 165.365 93.910 173.350 ;
        RECT 94.910 172.815 96.790 173.185 ;
        RECT 102.410 172.815 104.290 173.185 ;
        RECT 104.810 172.650 104.950 177.090 ;
        RECT 105.210 176.070 105.470 176.390 ;
        RECT 105.270 175.370 105.410 176.070 ;
        RECT 105.210 175.050 105.470 175.370 ;
        RECT 105.730 173.670 105.870 181.510 ;
        RECT 106.110 180.975 107.990 181.345 ;
        RECT 107.970 179.810 108.230 180.130 ;
        RECT 108.030 179.530 108.170 179.810 ;
        RECT 108.490 179.530 108.630 184.910 ;
        RECT 108.030 179.390 108.630 179.530 ;
        RECT 106.110 175.535 107.990 175.905 ;
        RECT 108.490 174.690 108.630 179.390 ;
        RECT 108.430 174.370 108.690 174.690 ;
        RECT 105.670 173.350 105.930 173.670 ;
        RECT 108.950 172.650 109.090 192.730 ;
        RECT 113.610 191.855 115.490 192.225 ;
        RECT 112.570 189.670 112.830 189.990 ;
        RECT 109.910 189.135 111.790 189.505 ;
        RECT 112.630 185.570 112.770 189.670 ;
        RECT 115.850 187.805 115.990 207.270 ;
        RECT 117.410 194.575 119.290 194.945 ;
        RECT 116.250 192.390 116.510 192.710 ;
        RECT 116.310 188.290 116.450 192.390 ;
        RECT 117.410 189.135 119.290 189.505 ;
        RECT 116.250 187.970 116.510 188.290 ;
        RECT 115.780 187.435 116.060 187.805 ;
        RECT 113.610 186.415 115.490 186.785 ;
        RECT 112.570 185.250 112.830 185.570 ;
        RECT 112.570 184.570 112.830 184.890 ;
        RECT 109.910 183.695 111.790 184.065 ;
        RECT 112.630 182.850 112.770 184.570 ;
        RECT 112.570 182.530 112.830 182.850 ;
        RECT 113.610 180.975 115.490 181.345 ;
        RECT 109.910 178.255 111.790 178.625 ;
        RECT 116.310 177.410 116.450 187.970 ;
        RECT 119.930 185.250 120.190 185.570 ;
        RECT 119.990 184.405 120.130 185.250 ;
        RECT 117.410 183.695 119.290 184.065 ;
        RECT 119.920 184.035 120.200 184.405 ;
        RECT 117.410 178.255 119.290 178.625 ;
        RECT 116.250 177.090 116.510 177.410 ;
        RECT 113.610 175.535 115.490 175.905 ;
        RECT 109.910 172.815 111.790 173.185 ;
        RECT 104.750 172.330 105.010 172.650 ;
        RECT 108.890 172.330 109.150 172.650 ;
        RECT 113.020 172.475 113.300 172.845 ;
        RECT 117.410 172.815 119.290 173.185 ;
        RECT 113.090 171.630 113.230 172.475 ;
        RECT 105.210 171.310 105.470 171.630 ;
        RECT 113.030 171.310 113.290 171.630 ;
        RECT 98.610 170.095 100.490 170.465 ;
        RECT 93.700 164.995 93.980 165.365 ;
        RECT 105.270 163.400 105.410 171.310 ;
        RECT 106.110 170.095 107.990 170.465 ;
        RECT 113.610 170.095 115.490 170.465 ;
        RECT 105.200 159.400 105.480 163.400 ;
        RECT 47.700 155.450 48.400 157.050 ;
        RECT 61.200 155.450 62.000 157.050 ;
        RECT 75.000 155.450 75.800 157.050 ;
        RECT 88.700 155.450 89.500 157.050 ;
        RECT 105.200 156.350 105.500 159.400 ;
        RECT 104.700 155.450 105.500 156.350 ;
        RECT 47.950 152.750 51.660 152.770 ;
        RECT 47.930 152.545 51.660 152.750 ;
        RECT 55.055 152.750 58.830 152.770 ;
        RECT 47.930 152.490 51.695 152.545 ;
        RECT 47.950 152.470 51.695 152.490 ;
        RECT 49.740 152.285 51.695 152.470 ;
        RECT 49.770 152.270 51.660 152.285 ;
        RECT 52.835 151.845 53.835 152.565 ;
        RECT 55.055 152.550 58.865 152.750 ;
        RECT 61.480 152.725 65.190 152.745 ;
        RECT 55.025 152.485 58.865 152.550 ;
        RECT 61.460 152.520 65.190 152.725 ;
        RECT 68.585 152.725 72.360 152.745 ;
        RECT 75.285 152.725 78.995 152.745 ;
        RECT 55.025 152.470 58.830 152.485 ;
        RECT 55.025 152.290 56.975 152.470 ;
        RECT 61.460 152.465 65.225 152.520 ;
        RECT 61.480 152.445 65.225 152.465 ;
        RECT 55.055 152.270 56.945 152.290 ;
        RECT 63.270 152.260 65.225 152.445 ;
        RECT 63.300 152.245 65.190 152.260 ;
        RECT 52.800 151.585 53.860 151.845 ;
        RECT 66.365 151.820 67.365 152.540 ;
        RECT 68.585 152.525 72.395 152.725 ;
        RECT 68.555 152.460 72.395 152.525 ;
        RECT 75.265 152.520 78.995 152.725 ;
        RECT 82.390 152.725 86.165 152.745 ;
        RECT 88.975 152.725 92.685 152.745 ;
        RECT 75.265 152.465 79.030 152.520 ;
        RECT 68.555 152.445 72.360 152.460 ;
        RECT 75.285 152.445 79.030 152.465 ;
        RECT 68.555 152.265 70.505 152.445 ;
        RECT 68.585 152.245 70.475 152.265 ;
        RECT 77.075 152.260 79.030 152.445 ;
        RECT 77.105 152.245 78.995 152.260 ;
        RECT 80.170 151.820 81.170 152.540 ;
        RECT 82.390 152.525 86.200 152.725 ;
        RECT 82.360 152.460 86.200 152.525 ;
        RECT 88.955 152.520 92.685 152.725 ;
        RECT 96.080 152.725 99.855 152.745 ;
        RECT 88.955 152.465 92.720 152.520 ;
        RECT 82.360 152.445 86.165 152.460 ;
        RECT 88.975 152.445 92.720 152.465 ;
        RECT 82.360 152.265 84.310 152.445 ;
        RECT 82.390 152.245 84.280 152.265 ;
        RECT 90.765 152.260 92.720 152.445 ;
        RECT 90.795 152.245 92.685 152.260 ;
        RECT 93.860 151.820 94.860 152.540 ;
        RECT 96.080 152.525 99.890 152.725 ;
        RECT 96.050 152.460 99.890 152.525 ;
        RECT 96.050 152.445 99.855 152.460 ;
        RECT 96.050 152.265 98.000 152.445 ;
        RECT 96.080 152.245 97.970 152.265 ;
        RECT 52.835 151.565 53.835 151.585 ;
        RECT 66.330 151.560 67.390 151.820 ;
        RECT 80.135 151.560 81.195 151.820 ;
        RECT 93.825 151.560 94.885 151.820 ;
        RECT 66.365 151.540 67.365 151.560 ;
        RECT 80.170 151.540 81.170 151.560 ;
        RECT 93.860 151.540 94.860 151.560 ;
        RECT 47.970 150.320 51.660 150.340 ;
        RECT 47.945 150.125 51.660 150.320 ;
        RECT 55.055 150.320 58.765 150.340 ;
        RECT 55.055 150.130 58.800 150.320 ;
        RECT 61.500 150.295 65.190 150.315 ;
        RECT 47.945 150.060 51.690 150.125 ;
        RECT 47.970 150.040 51.690 150.060 ;
        RECT 49.740 149.865 51.690 150.040 ;
        RECT 55.025 150.060 58.800 150.130 ;
        RECT 61.475 150.100 65.190 150.295 ;
        RECT 68.585 150.295 72.295 150.315 ;
        RECT 75.305 150.295 78.995 150.315 ;
        RECT 68.585 150.105 72.330 150.295 ;
        RECT 55.025 150.040 58.765 150.060 ;
        RECT 55.025 149.870 56.970 150.040 ;
        RECT 61.475 150.035 65.220 150.100 ;
        RECT 61.500 150.015 65.220 150.035 ;
        RECT 49.770 149.840 51.660 149.865 ;
        RECT 55.055 149.840 56.945 149.870 ;
        RECT 63.270 149.840 65.220 150.015 ;
        RECT 68.555 150.035 72.330 150.105 ;
        RECT 75.280 150.100 78.995 150.295 ;
        RECT 82.390 150.295 86.100 150.315 ;
        RECT 88.995 150.295 92.685 150.315 ;
        RECT 82.390 150.105 86.135 150.295 ;
        RECT 75.280 150.035 79.025 150.100 ;
        RECT 68.555 150.015 72.295 150.035 ;
        RECT 75.305 150.015 79.025 150.035 ;
        RECT 68.555 149.845 70.500 150.015 ;
        RECT 63.300 149.815 65.190 149.840 ;
        RECT 68.585 149.815 70.475 149.845 ;
        RECT 77.075 149.840 79.025 150.015 ;
        RECT 82.360 150.035 86.135 150.105 ;
        RECT 88.970 150.100 92.685 150.295 ;
        RECT 96.080 150.295 99.790 150.315 ;
        RECT 96.080 150.105 99.825 150.295 ;
        RECT 88.970 150.035 92.715 150.100 ;
        RECT 82.360 150.015 86.100 150.035 ;
        RECT 88.995 150.015 92.715 150.035 ;
        RECT 82.360 149.845 84.305 150.015 ;
        RECT 77.105 149.815 78.995 149.840 ;
        RECT 82.390 149.815 84.280 149.845 ;
        RECT 90.765 149.840 92.715 150.015 ;
        RECT 96.050 150.035 99.825 150.105 ;
        RECT 96.050 150.015 99.790 150.035 ;
        RECT 96.050 149.845 97.995 150.015 ;
        RECT 90.795 149.815 92.685 149.840 ;
        RECT 96.080 149.815 97.970 149.845 ;
        RECT 52.860 149.270 53.260 149.275 ;
        RECT 49.680 149.010 56.975 149.270 ;
        RECT 66.390 149.245 66.790 149.250 ;
        RECT 80.195 149.245 80.595 149.250 ;
        RECT 93.885 149.245 94.285 149.250 ;
        RECT 47.930 148.480 48.590 148.485 ;
        RECT 47.930 148.225 51.690 148.480 ;
        RECT 47.980 148.220 51.690 148.225 ;
        RECT 52.860 147.690 53.260 149.010 ;
        RECT 63.210 148.985 70.505 149.245 ;
        RECT 77.015 148.985 84.310 149.245 ;
        RECT 90.705 148.985 98.000 149.245 ;
        RECT 55.040 148.220 58.810 148.480 ;
        RECT 61.460 148.455 62.120 148.460 ;
        RECT 61.460 148.200 65.220 148.455 ;
        RECT 61.510 148.195 65.220 148.200 ;
        RECT 49.745 147.430 56.965 147.690 ;
        RECT 66.390 147.665 66.790 148.985 ;
        RECT 75.265 148.455 75.925 148.460 ;
        RECT 68.570 148.195 72.340 148.455 ;
        RECT 75.265 148.200 79.025 148.455 ;
        RECT 75.315 148.195 79.025 148.200 ;
        RECT 80.195 147.665 80.595 148.985 ;
        RECT 88.955 148.455 89.615 148.460 ;
        RECT 82.375 148.195 86.145 148.455 ;
        RECT 88.955 148.200 92.715 148.455 ;
        RECT 89.005 148.195 92.715 148.200 ;
        RECT 93.885 147.665 94.285 148.985 ;
        RECT 96.065 148.195 99.835 148.455 ;
        RECT 52.860 146.110 53.260 147.430 ;
        RECT 63.275 147.405 70.495 147.665 ;
        RECT 77.080 147.405 84.300 147.665 ;
        RECT 90.770 147.405 97.990 147.665 ;
        RECT 55.025 146.640 58.810 146.900 ;
        RECT 52.855 145.850 56.965 146.110 ;
        RECT 66.390 146.085 66.790 147.405 ;
        RECT 68.555 146.615 72.340 146.875 ;
        RECT 80.195 146.085 80.595 147.405 ;
        RECT 82.360 146.615 86.145 146.875 ;
        RECT 93.885 146.085 94.285 147.405 ;
        RECT 96.050 146.615 99.835 146.875 ;
        RECT 52.855 145.110 53.855 145.850 ;
        RECT 66.385 145.825 70.495 146.085 ;
        RECT 80.190 145.825 84.300 146.085 ;
        RECT 93.880 145.825 97.990 146.085 ;
        RECT 52.900 139.600 53.800 145.110 ;
        RECT 66.385 145.085 67.385 145.825 ;
        RECT 80.190 145.085 81.190 145.825 ;
        RECT 93.880 145.085 94.880 145.825 ;
        RECT 58.300 141.550 59.100 143.950 ;
        RECT 66.500 140.700 67.300 145.085 ;
        RECT 71.800 141.550 72.600 143.950 ;
        RECT 80.300 140.700 81.100 145.085 ;
        RECT 82.400 141.550 83.200 143.950 ;
        RECT 85.600 141.550 86.400 143.950 ;
        RECT 66.500 140.100 72.200 140.700 ;
        RECT 52.900 139.100 70.200 139.600 ;
        RECT 69.400 138.265 70.200 139.100 ;
        RECT 71.400 138.265 72.200 140.100 ;
        RECT 73.500 140.100 81.100 140.700 ;
        RECT 73.500 138.265 74.200 140.100 ;
        RECT 94.000 139.600 94.800 145.085 ;
        RECT 99.300 141.550 100.100 143.950 ;
        RECT 75.400 139.100 94.800 139.600 ;
        RECT 75.400 138.265 76.200 139.100 ;
        RECT 69.285 137.265 70.285 138.265 ;
        RECT 71.295 137.265 72.295 138.265 ;
        RECT 73.305 137.265 74.305 138.265 ;
        RECT 75.315 137.265 76.315 138.265 ;
        RECT 69.285 134.190 69.545 137.265 ;
        RECT 71.295 133.790 71.555 137.265 ;
        RECT 73.305 135.790 73.570 137.265 ;
        RECT 73.305 133.790 73.565 135.790 ;
        RECT 75.315 133.990 75.575 137.265 ;
        RECT 100.550 134.275 100.830 134.310 ;
        RECT 99.760 134.270 100.850 134.275 ;
        RECT 87.565 133.590 90.090 133.605 ;
        RECT 85.840 132.425 90.090 133.590 ;
        RECT 99.250 132.935 100.850 134.270 ;
        RECT 112.755 133.585 113.805 133.615 ;
        RECT 85.840 132.405 88.005 132.425 ;
        RECT 85.845 130.485 87.015 132.405 ;
        RECT 87.670 132.390 87.970 132.405 ;
        RECT 85.840 130.170 87.020 130.485 ;
        RECT 99.250 130.170 100.210 132.935 ;
        RECT 100.550 132.895 100.830 132.935 ;
        RECT 101.125 131.670 102.965 131.710 ;
        RECT 104.700 131.690 106.555 131.720 ;
        RECT 85.840 129.870 100.210 130.170 ;
        RECT 101.115 130.695 102.980 131.670 ;
        RECT 85.840 129.205 100.190 129.870 ;
        RECT 85.840 129.090 87.020 129.205 ;
        RECT 98.320 129.200 100.190 129.205 ;
        RECT 85.820 128.420 87.020 129.090 ;
        RECT 101.115 128.535 102.295 130.695 ;
        RECT 104.680 130.340 106.565 131.690 ;
        RECT 100.995 128.530 102.295 128.535 ;
        RECT 85.830 128.330 87.020 128.420 ;
        RECT 85.840 126.875 87.020 128.330 ;
        RECT 99.995 127.695 102.295 128.530 ;
        RECT 105.460 129.740 106.565 130.340 ;
        RECT 112.715 130.100 113.885 133.585 ;
        RECT 105.460 128.755 110.620 129.740 ;
        RECT 112.715 129.300 118.700 130.100 ;
        RECT 99.175 127.005 99.440 127.025 ;
        RECT 99.995 127.005 101.085 127.695 ;
        RECT 87.720 126.875 88.000 126.900 ;
        RECT 85.840 126.495 88.005 126.875 ;
        RECT 85.835 125.695 88.005 126.495 ;
        RECT 99.165 126.590 101.085 127.005 ;
        RECT 104.895 127.010 105.190 127.045 ;
        RECT 105.460 127.010 106.565 128.755 ;
        RECT 99.165 125.820 101.075 126.590 ;
        RECT 104.895 125.920 106.565 127.010 ;
        RECT 104.895 125.885 105.190 125.920 ;
        RECT 99.175 125.805 99.440 125.820 ;
        RECT 100.860 125.815 101.075 125.820 ;
        RECT 112.715 125.720 113.885 129.300 ;
        RECT 112.715 125.695 113.845 125.720 ;
        RECT 86.045 125.690 88.005 125.695 ;
        RECT 87.720 125.640 88.000 125.690 ;
        RECT 102.600 125.525 102.870 125.555 ;
        RECT 107.070 125.525 107.335 125.555 ;
        RECT 96.880 125.485 97.150 125.520 ;
        RECT 101.320 125.485 101.630 125.525 ;
        RECT 102.595 125.520 107.350 125.525 ;
        RECT 94.775 125.470 96.020 125.475 ;
        RECT 96.880 125.470 101.650 125.485 ;
        RECT 94.775 124.585 101.650 125.470 ;
        RECT 67.290 123.995 67.550 124.035 ;
        RECT 69.240 123.995 69.500 124.035 ;
        RECT 67.280 122.035 69.515 123.995 ;
        RECT 67.280 122.025 69.545 122.035 ;
        RECT 67.290 121.985 67.550 122.025 ;
        RECT 69.240 121.985 69.545 122.025 ;
        RECT 69.285 118.170 69.545 121.985 ;
        RECT 71.295 120.130 71.555 124.045 ;
        RECT 73.305 123.945 73.565 124.045 ;
        RECT 70.335 118.260 71.555 120.130 ;
        RECT 67.100 111.150 67.700 116.950 ;
        RECT 69.285 113.380 69.545 113.425 ;
        RECT 70.335 113.380 70.535 118.260 ;
        RECT 71.295 118.170 71.555 118.260 ;
        RECT 72.330 122.075 73.565 123.945 ;
        RECT 69.285 111.510 70.535 113.380 ;
        RECT 71.295 113.345 71.555 113.425 ;
        RECT 72.330 113.345 72.530 122.075 ;
        RECT 73.305 121.995 73.565 122.075 ;
        RECT 73.305 120.150 73.565 120.220 ;
        RECT 75.315 120.150 75.575 124.045 ;
        RECT 88.165 122.645 89.970 123.015 ;
        RECT 73.305 120.000 75.575 120.150 ;
        RECT 88.315 120.000 89.780 122.645 ;
        RECT 91.615 122.635 93.420 123.005 ;
        RECT 73.305 119.200 89.780 120.000 ;
        RECT 73.305 119.150 75.575 119.200 ;
        RECT 73.305 118.170 73.565 119.150 ;
        RECT 88.315 119.010 89.780 119.200 ;
        RECT 91.765 118.985 93.230 122.635 ;
        RECT 94.775 121.815 96.020 124.585 ;
        RECT 96.880 124.560 101.650 124.585 ;
        RECT 102.595 124.580 109.310 125.520 ;
        RECT 102.595 124.570 107.350 124.580 ;
        RECT 96.880 124.530 97.150 124.560 ;
        RECT 101.320 124.520 101.630 124.560 ;
        RECT 102.600 124.535 102.870 124.570 ;
        RECT 107.070 124.530 107.335 124.570 ;
        RECT 103.560 124.290 103.855 124.295 ;
        RECT 106.030 124.290 106.290 124.295 ;
        RECT 103.485 124.280 106.440 124.290 ;
        RECT 98.140 124.275 98.440 124.280 ;
        RECT 100.200 124.275 106.440 124.280 ;
        RECT 98.050 123.315 106.440 124.275 ;
        RECT 98.050 123.305 100.610 123.315 ;
        RECT 108.290 121.880 109.310 124.580 ;
        RECT 108.350 121.870 109.240 121.880 ;
        RECT 94.805 121.800 95.950 121.815 ;
        RECT 118.000 120.400 118.700 129.300 ;
        RECT 122.665 122.635 123.020 122.660 ;
        RECT 120.020 121.890 120.280 121.925 ;
        RECT 119.970 120.590 120.280 121.890 ;
        RECT 121.395 121.870 121.695 121.910 ;
        RECT 119.290 120.400 120.300 120.590 ;
        RECT 118.000 119.700 120.300 120.400 ;
        RECT 121.385 119.930 121.980 121.870 ;
        RECT 122.635 120.860 123.050 122.635 ;
        RECT 122.635 120.825 123.225 120.860 ;
        RECT 124.360 120.825 124.630 120.860 ;
        RECT 122.635 119.935 123.240 120.825 ;
        RECT 124.345 119.935 124.955 120.825 ;
        RECT 121.395 119.890 121.980 119.930 ;
        RECT 122.965 119.905 123.225 119.935 ;
        RECT 124.360 119.900 124.955 119.935 ;
        RECT 119.290 119.590 120.300 119.700 ;
        RECT 119.955 118.400 120.955 118.595 ;
        RECT 116.300 117.800 120.955 118.400 ;
        RECT 119.955 117.595 120.955 117.800 ;
        RECT 121.625 118.320 121.980 119.890 ;
        RECT 124.550 118.595 124.955 119.900 ;
        RECT 122.915 118.320 123.195 118.345 ;
        RECT 121.625 117.920 123.220 118.320 ;
        RECT 119.285 116.600 120.295 116.725 ;
        RECT 117.500 115.800 120.295 116.600 ;
        RECT 121.625 116.415 121.980 117.920 ;
        RECT 122.915 117.900 123.195 117.920 ;
        RECT 124.545 117.595 125.555 118.595 ;
        RECT 121.400 116.375 121.980 116.415 ;
        RECT 73.305 113.345 73.565 113.425 ;
        RECT 69.285 111.375 69.545 111.510 ;
        RECT 71.295 111.460 73.565 113.345 ;
        RECT 71.295 111.375 71.555 111.460 ;
        RECT 73.305 111.375 73.565 111.460 ;
        RECT 46.600 108.050 48.400 108.950 ;
        RECT 82.925 102.645 83.185 113.370 ;
        RECT 89.805 111.415 90.065 111.440 ;
        RECT 93.665 111.425 93.925 111.455 ;
        RECT 89.495 109.460 90.095 111.415 ;
        RECT 93.635 109.460 94.235 111.425 ;
        RECT 89.495 109.435 90.065 109.460 ;
        RECT 93.665 109.440 94.235 109.460 ;
        RECT 84.845 108.190 85.115 108.240 ;
        RECT 89.495 108.190 89.895 109.435 ;
        RECT 90.245 108.190 90.560 108.240 ;
        RECT 93.160 108.195 93.490 108.245 ;
        RECT 93.835 108.195 94.235 109.440 ;
        RECT 98.630 108.195 98.900 108.245 ;
        RECT 84.830 107.930 90.580 108.190 ;
        RECT 84.845 107.880 85.115 107.930 ;
        RECT 86.595 107.790 90.580 107.930 ;
        RECT 93.145 107.935 98.915 108.195 ;
        RECT 93.145 107.795 97.135 107.935 ;
        RECT 98.630 107.885 98.900 107.935 ;
        RECT 86.595 104.570 86.895 107.790 ;
        RECT 88.505 106.075 89.505 107.075 ;
        RECT 93.520 106.075 94.520 107.075 ;
        RECT 89.035 106.060 89.475 106.075 ;
        RECT 94.060 106.065 94.475 106.075 ;
        RECT 96.835 104.570 97.135 107.795 ;
        RECT 86.595 104.550 87.065 104.570 ;
        RECT 86.600 102.650 87.100 104.550 ;
        RECT 96.665 104.545 97.135 104.570 ;
        RECT 96.635 102.655 97.135 104.545 ;
        RECT 86.805 102.640 87.065 102.650 ;
        RECT 96.665 102.635 96.925 102.655 ;
        RECT 100.555 102.630 100.815 113.380 ;
        RECT 105.370 110.370 105.630 110.410 ;
        RECT 105.345 109.980 105.845 110.370 ;
        RECT 105.370 109.940 105.845 109.980 ;
        RECT 105.545 108.745 105.845 109.940 ;
        RECT 105.540 108.700 106.540 108.745 ;
        RECT 117.500 108.700 118.400 115.800 ;
        RECT 119.285 115.725 120.295 115.800 ;
        RECT 119.970 114.440 120.280 115.725 ;
        RECT 120.020 114.425 120.280 114.440 ;
        RECT 121.385 114.430 121.980 116.375 ;
        RECT 122.960 116.370 123.220 116.405 ;
        RECT 124.550 116.395 124.955 117.595 ;
        RECT 124.365 116.375 124.955 116.395 ;
        RECT 122.640 115.480 123.235 116.370 ;
        RECT 124.345 115.480 124.955 116.375 ;
        RECT 122.640 115.445 123.220 115.480 ;
        RECT 124.365 115.465 124.635 115.480 ;
        RECT 121.400 114.395 121.700 114.430 ;
        RECT 122.640 113.850 123.055 115.445 ;
        RECT 122.670 113.830 123.030 113.850 ;
        RECT 105.540 107.800 118.400 108.700 ;
        RECT 105.540 107.745 106.540 107.800 ;
        RECT 105.545 106.575 105.845 107.745 ;
        RECT 105.380 106.540 105.845 106.575 ;
        RECT 105.345 105.690 105.845 106.540 ;
        RECT 105.380 105.655 105.640 105.690 ;
        RECT 80.100 100.250 89.700 101.150 ;
      LAYER met3 ;
        RECT 68.100 194.000 68.700 220.600 ;
        RECT 72.700 218.600 73.900 219.200 ;
        RECT 78.300 217.300 79.500 217.900 ;
        RECT 88.200 203.560 88.800 214.000 ;
        RECT 140.850 213.075 141.450 213.625 ;
        RECT 143.650 210.475 144.250 211.025 ;
        RECT 85.330 203.410 89.330 203.560 ;
        RECT 92.295 203.410 92.625 203.425 ;
        RECT 85.330 203.110 92.625 203.410 ;
        RECT 85.330 202.960 89.330 203.110 ;
        RECT 92.295 203.095 92.625 203.110 ;
        RECT 98.560 197.315 100.540 197.645 ;
        RECT 106.060 197.315 108.040 197.645 ;
        RECT 113.560 197.315 115.540 197.645 ;
        RECT 94.860 194.595 96.840 194.925 ;
        RECT 102.360 194.595 104.340 194.925 ;
        RECT 109.860 194.595 111.840 194.925 ;
        RECT 117.360 194.595 119.340 194.925 ;
        RECT 85.330 194.000 89.330 194.040 ;
        RECT 53.000 193.890 89.330 194.000 ;
        RECT 93.675 193.890 94.005 193.905 ;
        RECT 53.000 193.590 94.005 193.890 ;
        RECT 53.000 193.440 89.330 193.590 ;
        RECT 93.675 193.575 94.005 193.590 ;
        RECT 53.000 193.400 85.400 193.440 ;
        RECT 47.650 155.475 48.450 157.025 ;
        RECT 53.000 151.700 53.600 193.400 ;
        RECT 98.560 191.875 100.540 192.205 ;
        RECT 106.060 191.875 108.040 192.205 ;
        RECT 113.560 191.875 115.540 192.205 ;
        RECT 94.860 189.155 96.840 189.485 ;
        RECT 102.360 189.155 104.340 189.485 ;
        RECT 109.860 189.155 111.840 189.485 ;
        RECT 117.360 189.155 119.340 189.485 ;
        RECT 115.755 187.780 116.085 187.785 ;
        RECT 115.755 187.770 116.340 187.780 ;
        RECT 115.530 187.470 116.340 187.770 ;
        RECT 115.755 187.460 116.340 187.470 ;
        RECT 115.755 187.455 116.085 187.460 ;
        RECT 98.560 186.435 100.540 186.765 ;
        RECT 106.060 186.435 108.040 186.765 ;
        RECT 113.560 186.435 115.540 186.765 ;
        RECT 72.700 184.500 73.300 185.100 ;
        RECT 89.535 185.050 89.865 185.065 ;
        RECT 89.320 184.735 89.865 185.050 ;
        RECT 89.320 184.520 89.620 184.735 ;
        RECT 125.200 184.520 127.100 184.600 ;
        RECT 85.330 184.500 89.620 184.520 ;
        RECT 66.500 184.070 89.620 184.500 ;
        RECT 119.895 184.370 120.225 184.385 ;
        RECT 121.965 184.370 127.100 184.520 ;
        RECT 119.895 184.070 127.100 184.370 ;
        RECT 66.500 183.920 89.330 184.070 ;
        RECT 119.895 184.055 120.225 184.070 ;
        RECT 66.500 183.900 85.600 183.920 ;
        RECT 61.150 155.475 62.050 157.025 ;
        RECT 66.500 151.700 67.200 183.900 ;
        RECT 94.860 183.715 96.840 184.045 ;
        RECT 102.360 183.715 104.340 184.045 ;
        RECT 109.860 183.715 111.840 184.045 ;
        RECT 117.360 183.715 119.340 184.045 ;
        RECT 121.965 183.920 127.100 184.070 ;
        RECT 125.200 183.800 127.100 183.920 ;
        RECT 98.560 180.995 100.540 181.325 ;
        RECT 106.060 180.995 108.040 181.325 ;
        RECT 113.560 180.995 115.540 181.325 ;
        RECT 94.860 178.275 96.840 178.605 ;
        RECT 102.360 178.275 104.340 178.605 ;
        RECT 109.860 178.275 111.840 178.605 ;
        RECT 117.360 178.275 119.340 178.605 ;
        RECT 98.560 175.555 100.540 175.885 ;
        RECT 106.060 175.555 108.040 175.885 ;
        RECT 113.560 175.555 115.540 175.885 ;
        RECT 77.700 174.850 89.330 175.000 ;
        RECT 77.700 174.400 89.620 174.850 ;
        RECT 74.950 155.475 75.850 157.025 ;
        RECT 80.300 151.800 81.000 174.400 ;
        RECT 89.320 174.185 89.620 174.400 ;
        RECT 89.320 173.870 89.865 174.185 ;
        RECT 89.535 173.855 89.865 173.870 ;
        RECT 94.860 172.835 96.840 173.165 ;
        RECT 102.360 172.835 104.340 173.165 ;
        RECT 109.860 172.835 111.840 173.165 ;
        RECT 117.360 172.835 119.340 173.165 ;
        RECT 112.995 172.810 113.325 172.825 ;
        RECT 115.960 172.810 116.340 172.820 ;
        RECT 112.995 172.510 116.340 172.810 ;
        RECT 112.995 172.495 113.325 172.510 ;
        RECT 115.960 172.500 116.340 172.510 ;
        RECT 98.560 170.115 100.540 170.445 ;
        RECT 106.060 170.115 108.040 170.445 ;
        RECT 113.560 170.115 115.540 170.445 ;
        RECT 87.600 165.480 88.500 165.500 ;
        RECT 85.330 165.330 89.330 165.480 ;
        RECT 93.675 165.330 94.005 165.345 ;
        RECT 85.330 165.030 94.005 165.330 ;
        RECT 85.330 164.880 89.330 165.030 ;
        RECT 93.675 165.015 94.005 165.030 ;
        RECT 87.600 162.900 88.500 164.880 ;
        RECT 87.600 162.400 94.600 162.900 ;
        RECT 94.000 158.000 94.600 162.400 ;
        RECT 94.000 157.500 116.900 158.000 ;
        RECT 88.650 155.475 89.550 157.025 ;
        RECT 94.000 151.700 94.700 157.500 ;
        RECT 104.650 155.475 105.550 156.325 ;
        RECT 1.400 144.000 45.900 144.100 ;
        RECT 1.400 141.500 100.200 144.000 ;
        RECT 1.400 141.400 45.800 141.500 ;
        RECT 46.500 108.000 48.500 141.500 ;
        RECT 67.050 111.175 67.750 116.925 ;
        RECT 87.500 107.000 88.200 120.000 ;
        RECT 92.100 119.300 109.400 120.200 ;
        RECT 87.500 106.200 89.400 107.000 ;
        RECT 80.050 100.275 89.750 101.125 ;
        RECT 93.700 94.200 94.400 106.900 ;
        RECT 108.700 94.200 109.400 119.300 ;
        RECT 116.300 117.800 116.900 157.500 ;
        RECT 126.300 118.500 127.100 183.800 ;
        RECT 124.600 117.700 127.100 118.500 ;
        RECT 93.700 93.200 152.700 94.200 ;
      LAYER met4 ;
        RECT 83.000 224.760 83.110 224.900 ;
        RECT 83.410 224.760 83.500 224.900 ;
        RECT 83.000 220.600 83.500 224.760 ;
        RECT 68.100 220.000 83.500 220.600 ;
        RECT 85.800 224.760 85.870 224.900 ;
        RECT 86.170 224.760 86.200 224.900 ;
        RECT 85.800 219.200 86.200 224.760 ;
        RECT 73.300 218.600 86.200 219.200 ;
        RECT 88.600 224.760 88.630 224.900 ;
        RECT 88.930 224.760 89.000 224.900 ;
        RECT 88.600 217.900 89.000 224.760 ;
        RECT 78.900 217.300 89.000 217.900 ;
        RECT 91.300 224.760 91.390 224.800 ;
        RECT 91.690 224.760 91.800 224.800 ;
        RECT 91.300 215.900 91.800 224.760 ;
        RECT 83.100 215.300 91.800 215.900 ;
        RECT 94.100 224.760 94.150 224.800 ;
        RECT 94.450 224.760 94.500 224.800 ;
        RECT 83.100 165.500 83.600 215.300 ;
        RECT 88.200 213.900 89.000 214.000 ;
        RECT 94.100 213.900 94.500 224.760 ;
        RECT 88.200 213.400 94.500 213.900 ;
        RECT 141.000 224.760 141.070 224.900 ;
        RECT 141.370 224.760 141.400 224.900 ;
        RECT 141.000 213.700 141.400 224.760 ;
        RECT 143.700 224.760 143.830 224.900 ;
        RECT 144.130 224.760 144.200 224.900 ;
        RECT 140.800 213.000 141.500 213.700 ;
        RECT 143.700 211.100 144.200 224.760 ;
        RECT 143.600 210.400 144.300 211.100 ;
        RECT 94.850 170.040 96.850 197.720 ;
        RECT 98.550 170.040 100.550 197.720 ;
        RECT 102.350 170.040 104.350 197.720 ;
        RECT 106.050 170.040 108.050 197.720 ;
        RECT 109.850 170.040 111.850 197.720 ;
        RECT 113.550 170.040 115.550 197.720 ;
        RECT 115.985 187.455 116.315 187.785 ;
        RECT 116.000 172.825 116.300 187.455 ;
        RECT 115.985 172.495 116.315 172.825 ;
        RECT 117.350 170.040 119.350 197.720 ;
        RECT 83.100 164.900 85.900 165.500 ;
        RECT 6.000 156.400 89.800 157.100 ;
        RECT 6.000 155.400 105.700 156.400 ;
        RECT 66.900 101.200 67.800 117.000 ;
        RECT 6.000 100.200 90.100 101.200 ;
        RECT 151.775 1.000 152.765 94.285 ;
        RECT 151.775 0.925 151.810 1.000 ;
        RECT 152.710 0.925 152.765 1.000 ;
      LAYER met5 ;
        RECT 90.610 192.980 120.530 194.980 ;
        RECT 90.610 189.280 120.530 191.280 ;
        RECT 90.610 185.480 120.530 187.480 ;
        RECT 90.610 181.780 120.530 183.780 ;
        RECT 90.610 177.980 120.530 179.980 ;
        RECT 90.610 174.280 120.530 176.280 ;
  END
END tt_um_4Bit_SAR_ADC
END LIBRARY

